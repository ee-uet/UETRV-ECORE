VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Motor_Top
  CLASS BLOCK ;
  FOREIGN Motor_Top ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 496.000 17.850 500.000 ;
    END
  END clock
  PIN io_ba_match
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 453.600 4.000 454.200 ;
    END
  END io_ba_match
  PIN io_motor_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END io_motor_irq
  PIN io_pwm_high
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 22.480 500.000 23.080 ;
    END
  END io_pwm_high
  PIN io_pwm_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 67.360 500.000 67.960 ;
    END
  END io_pwm_low
  PIN io_qei_ch_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END io_qei_ch_a
  PIN io_qei_ch_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END io_qei_ch_b
  PIN io_wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END io_wbs_ack_o
  PIN io_wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 496.000 89.150 500.000 ;
    END
  END io_wbs_data_o[0]
  PIN io_wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 204.040 500.000 204.640 ;
    END
  END io_wbs_data_o[10]
  PIN io_wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END io_wbs_data_o[11]
  PIN io_wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 496.000 267.630 500.000 ;
    END
  END io_wbs_data_o[12]
  PIN io_wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 496.000 303.510 500.000 ;
    END
  END io_wbs_data_o[13]
  PIN io_wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 249.600 500.000 250.200 ;
    END
  END io_wbs_data_o[14]
  PIN io_wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 496.000 338.930 500.000 ;
    END
  END io_wbs_data_o[15]
  PIN io_wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END io_wbs_data_o[16]
  PIN io_wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 496.000 374.810 500.000 ;
    END
  END io_wbs_data_o[17]
  PIN io_wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 294.480 500.000 295.080 ;
    END
  END io_wbs_data_o[18]
  PIN io_wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 340.040 500.000 340.640 ;
    END
  END io_wbs_data_o[19]
  PIN io_wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 496.000 124.570 500.000 ;
    END
  END io_wbs_data_o[1]
  PIN io_wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 496.000 410.690 500.000 ;
    END
  END io_wbs_data_o[20]
  PIN io_wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 496.000 446.110 500.000 ;
    END
  END io_wbs_data_o[21]
  PIN io_wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 496.000 481.990 500.000 ;
    END
  END io_wbs_data_o[22]
  PIN io_wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END io_wbs_data_o[23]
  PIN io_wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END io_wbs_data_o[24]
  PIN io_wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 385.600 500.000 386.200 ;
    END
  END io_wbs_data_o[25]
  PIN io_wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END io_wbs_data_o[26]
  PIN io_wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 431.160 500.000 431.760 ;
    END
  END io_wbs_data_o[27]
  PIN io_wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 476.720 500.000 477.320 ;
    END
  END io_wbs_data_o[28]
  PIN io_wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END io_wbs_data_o[29]
  PIN io_wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.760 4.000 462.360 ;
    END
  END io_wbs_data_o[2]
  PIN io_wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END io_wbs_data_o[30]
  PIN io_wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END io_wbs_data_o[31]
  PIN io_wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 496.000 160.450 500.000 ;
    END
  END io_wbs_data_o[3]
  PIN io_wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 496.000 196.330 500.000 ;
    END
  END io_wbs_data_o[4]
  PIN io_wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 112.920 500.000 113.520 ;
    END
  END io_wbs_data_o[5]
  PIN io_wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END io_wbs_data_o[6]
  PIN io_wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END io_wbs_data_o[7]
  PIN io_wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 496.000 231.750 500.000 ;
    END
  END io_wbs_data_o[8]
  PIN io_wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 158.480 500.000 159.080 ;
    END
  END io_wbs_data_o[9]
  PIN io_wbs_m2s_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END io_wbs_m2s_addr[0]
  PIN io_wbs_m2s_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END io_wbs_m2s_addr[10]
  PIN io_wbs_m2s_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END io_wbs_m2s_addr[11]
  PIN io_wbs_m2s_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 4.000 254.280 ;
    END
  END io_wbs_m2s_addr[12]
  PIN io_wbs_m2s_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END io_wbs_m2s_addr[13]
  PIN io_wbs_m2s_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END io_wbs_m2s_addr[14]
  PIN io_wbs_m2s_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.000 4.000 304.600 ;
    END
  END io_wbs_m2s_addr[15]
  PIN io_wbs_m2s_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END io_wbs_m2s_addr[1]
  PIN io_wbs_m2s_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END io_wbs_m2s_addr[2]
  PIN io_wbs_m2s_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END io_wbs_m2s_addr[3]
  PIN io_wbs_m2s_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END io_wbs_m2s_addr[4]
  PIN io_wbs_m2s_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END io_wbs_m2s_addr[5]
  PIN io_wbs_m2s_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END io_wbs_m2s_addr[6]
  PIN io_wbs_m2s_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END io_wbs_m2s_addr[7]
  PIN io_wbs_m2s_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END io_wbs_m2s_addr[8]
  PIN io_wbs_m2s_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END io_wbs_m2s_addr[9]
  PIN io_wbs_m2s_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END io_wbs_m2s_data[0]
  PIN io_wbs_m2s_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END io_wbs_m2s_data[10]
  PIN io_wbs_m2s_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END io_wbs_m2s_data[11]
  PIN io_wbs_m2s_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END io_wbs_m2s_data[12]
  PIN io_wbs_m2s_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END io_wbs_m2s_data[13]
  PIN io_wbs_m2s_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END io_wbs_m2s_data[14]
  PIN io_wbs_m2s_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END io_wbs_m2s_data[15]
  PIN io_wbs_m2s_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END io_wbs_m2s_data[16]
  PIN io_wbs_m2s_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END io_wbs_m2s_data[17]
  PIN io_wbs_m2s_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END io_wbs_m2s_data[18]
  PIN io_wbs_m2s_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END io_wbs_m2s_data[19]
  PIN io_wbs_m2s_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END io_wbs_m2s_data[1]
  PIN io_wbs_m2s_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END io_wbs_m2s_data[20]
  PIN io_wbs_m2s_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END io_wbs_m2s_data[21]
  PIN io_wbs_m2s_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END io_wbs_m2s_data[22]
  PIN io_wbs_m2s_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END io_wbs_m2s_data[23]
  PIN io_wbs_m2s_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END io_wbs_m2s_data[24]
  PIN io_wbs_m2s_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END io_wbs_m2s_data[25]
  PIN io_wbs_m2s_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END io_wbs_m2s_data[26]
  PIN io_wbs_m2s_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END io_wbs_m2s_data[27]
  PIN io_wbs_m2s_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END io_wbs_m2s_data[28]
  PIN io_wbs_m2s_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END io_wbs_m2s_data[29]
  PIN io_wbs_m2s_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END io_wbs_m2s_data[2]
  PIN io_wbs_m2s_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.280 4.000 437.880 ;
    END
  END io_wbs_m2s_data[30]
  PIN io_wbs_m2s_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END io_wbs_m2s_data[31]
  PIN io_wbs_m2s_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END io_wbs_m2s_data[3]
  PIN io_wbs_m2s_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END io_wbs_m2s_data[4]
  PIN io_wbs_m2s_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END io_wbs_m2s_data[5]
  PIN io_wbs_m2s_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END io_wbs_m2s_data[6]
  PIN io_wbs_m2s_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END io_wbs_m2s_data[7]
  PIN io_wbs_m2s_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END io_wbs_m2s_data[8]
  PIN io_wbs_m2s_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END io_wbs_m2s_data[9]
  PIN io_wbs_m2s_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END io_wbs_m2s_sel[0]
  PIN io_wbs_m2s_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END io_wbs_m2s_sel[1]
  PIN io_wbs_m2s_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END io_wbs_m2s_sel[2]
  PIN io_wbs_m2s_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END io_wbs_m2s_sel[3]
  PIN io_wbs_m2s_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END io_wbs_m2s_stb
  PIN io_wbs_m2s_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END io_wbs_m2s_we
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 496.000 53.270 500.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 5.520 10.640 494.040 487.120 ;
      LAYER met2 ;
        RECT 6.990 495.720 17.290 496.810 ;
        RECT 18.130 495.720 52.710 496.810 ;
        RECT 53.550 495.720 88.590 496.810 ;
        RECT 89.430 495.720 124.010 496.810 ;
        RECT 124.850 495.720 159.890 496.810 ;
        RECT 160.730 495.720 195.770 496.810 ;
        RECT 196.610 495.720 231.190 496.810 ;
        RECT 232.030 495.720 267.070 496.810 ;
        RECT 267.910 495.720 302.950 496.810 ;
        RECT 303.790 495.720 338.370 496.810 ;
        RECT 339.210 495.720 374.250 496.810 ;
        RECT 375.090 495.720 410.130 496.810 ;
        RECT 410.970 495.720 445.550 496.810 ;
        RECT 446.390 495.720 481.430 496.810 ;
        RECT 482.270 495.720 491.190 496.810 ;
        RECT 6.990 4.280 491.190 495.720 ;
        RECT 6.990 4.000 24.650 4.280 ;
        RECT 25.490 4.000 74.330 4.280 ;
        RECT 75.170 4.000 124.470 4.280 ;
        RECT 125.310 4.000 174.610 4.280 ;
        RECT 175.450 4.000 224.290 4.280 ;
        RECT 225.130 4.000 274.430 4.280 ;
        RECT 275.270 4.000 324.570 4.280 ;
        RECT 325.410 4.000 374.250 4.280 ;
        RECT 375.090 4.000 424.390 4.280 ;
        RECT 425.230 4.000 474.530 4.280 ;
        RECT 475.370 4.000 491.190 4.280 ;
      LAYER met3 ;
        RECT 4.400 494.680 496.000 495.545 ;
        RECT 4.000 487.920 496.000 494.680 ;
        RECT 4.400 486.520 496.000 487.920 ;
        RECT 4.000 479.760 496.000 486.520 ;
        RECT 4.400 478.360 496.000 479.760 ;
        RECT 4.000 477.720 496.000 478.360 ;
        RECT 4.000 476.320 495.600 477.720 ;
        RECT 4.000 471.600 496.000 476.320 ;
        RECT 4.400 470.200 496.000 471.600 ;
        RECT 4.000 462.760 496.000 470.200 ;
        RECT 4.400 461.360 496.000 462.760 ;
        RECT 4.000 454.600 496.000 461.360 ;
        RECT 4.400 453.200 496.000 454.600 ;
        RECT 4.000 446.440 496.000 453.200 ;
        RECT 4.400 445.040 496.000 446.440 ;
        RECT 4.000 438.280 496.000 445.040 ;
        RECT 4.400 436.880 496.000 438.280 ;
        RECT 4.000 432.160 496.000 436.880 ;
        RECT 4.000 430.760 495.600 432.160 ;
        RECT 4.000 429.440 496.000 430.760 ;
        RECT 4.400 428.040 496.000 429.440 ;
        RECT 4.000 421.280 496.000 428.040 ;
        RECT 4.400 419.880 496.000 421.280 ;
        RECT 4.000 413.120 496.000 419.880 ;
        RECT 4.400 411.720 496.000 413.120 ;
        RECT 4.000 404.960 496.000 411.720 ;
        RECT 4.400 403.560 496.000 404.960 ;
        RECT 4.000 396.120 496.000 403.560 ;
        RECT 4.400 394.720 496.000 396.120 ;
        RECT 4.000 387.960 496.000 394.720 ;
        RECT 4.400 386.600 496.000 387.960 ;
        RECT 4.400 386.560 495.600 386.600 ;
        RECT 4.000 385.200 495.600 386.560 ;
        RECT 4.000 379.800 496.000 385.200 ;
        RECT 4.400 378.400 496.000 379.800 ;
        RECT 4.000 371.640 496.000 378.400 ;
        RECT 4.400 370.240 496.000 371.640 ;
        RECT 4.000 362.800 496.000 370.240 ;
        RECT 4.400 361.400 496.000 362.800 ;
        RECT 4.000 354.640 496.000 361.400 ;
        RECT 4.400 353.240 496.000 354.640 ;
        RECT 4.000 346.480 496.000 353.240 ;
        RECT 4.400 345.080 496.000 346.480 ;
        RECT 4.000 341.040 496.000 345.080 ;
        RECT 4.000 339.640 495.600 341.040 ;
        RECT 4.000 338.320 496.000 339.640 ;
        RECT 4.400 336.920 496.000 338.320 ;
        RECT 4.000 329.480 496.000 336.920 ;
        RECT 4.400 328.080 496.000 329.480 ;
        RECT 4.000 321.320 496.000 328.080 ;
        RECT 4.400 319.920 496.000 321.320 ;
        RECT 4.000 313.160 496.000 319.920 ;
        RECT 4.400 311.760 496.000 313.160 ;
        RECT 4.000 305.000 496.000 311.760 ;
        RECT 4.400 303.600 496.000 305.000 ;
        RECT 4.000 296.160 496.000 303.600 ;
        RECT 4.400 295.480 496.000 296.160 ;
        RECT 4.400 294.760 495.600 295.480 ;
        RECT 4.000 294.080 495.600 294.760 ;
        RECT 4.000 288.000 496.000 294.080 ;
        RECT 4.400 286.600 496.000 288.000 ;
        RECT 4.000 279.840 496.000 286.600 ;
        RECT 4.400 278.440 496.000 279.840 ;
        RECT 4.000 271.680 496.000 278.440 ;
        RECT 4.400 270.280 496.000 271.680 ;
        RECT 4.000 262.840 496.000 270.280 ;
        RECT 4.400 261.440 496.000 262.840 ;
        RECT 4.000 254.680 496.000 261.440 ;
        RECT 4.400 253.280 496.000 254.680 ;
        RECT 4.000 250.600 496.000 253.280 ;
        RECT 4.000 249.200 495.600 250.600 ;
        RECT 4.000 246.520 496.000 249.200 ;
        RECT 4.400 245.120 496.000 246.520 ;
        RECT 4.000 238.360 496.000 245.120 ;
        RECT 4.400 236.960 496.000 238.360 ;
        RECT 4.000 229.520 496.000 236.960 ;
        RECT 4.400 228.120 496.000 229.520 ;
        RECT 4.000 221.360 496.000 228.120 ;
        RECT 4.400 219.960 496.000 221.360 ;
        RECT 4.000 213.200 496.000 219.960 ;
        RECT 4.400 211.800 496.000 213.200 ;
        RECT 4.000 205.040 496.000 211.800 ;
        RECT 4.400 203.640 495.600 205.040 ;
        RECT 4.000 196.200 496.000 203.640 ;
        RECT 4.400 194.800 496.000 196.200 ;
        RECT 4.000 188.040 496.000 194.800 ;
        RECT 4.400 186.640 496.000 188.040 ;
        RECT 4.000 179.880 496.000 186.640 ;
        RECT 4.400 178.480 496.000 179.880 ;
        RECT 4.000 171.720 496.000 178.480 ;
        RECT 4.400 170.320 496.000 171.720 ;
        RECT 4.000 162.880 496.000 170.320 ;
        RECT 4.400 161.480 496.000 162.880 ;
        RECT 4.000 159.480 496.000 161.480 ;
        RECT 4.000 158.080 495.600 159.480 ;
        RECT 4.000 154.720 496.000 158.080 ;
        RECT 4.400 153.320 496.000 154.720 ;
        RECT 4.000 146.560 496.000 153.320 ;
        RECT 4.400 145.160 496.000 146.560 ;
        RECT 4.000 138.400 496.000 145.160 ;
        RECT 4.400 137.000 496.000 138.400 ;
        RECT 4.000 129.560 496.000 137.000 ;
        RECT 4.400 128.160 496.000 129.560 ;
        RECT 4.000 121.400 496.000 128.160 ;
        RECT 4.400 120.000 496.000 121.400 ;
        RECT 4.000 113.920 496.000 120.000 ;
        RECT 4.000 113.240 495.600 113.920 ;
        RECT 4.400 112.520 495.600 113.240 ;
        RECT 4.400 111.840 496.000 112.520 ;
        RECT 4.000 105.080 496.000 111.840 ;
        RECT 4.400 103.680 496.000 105.080 ;
        RECT 4.000 96.240 496.000 103.680 ;
        RECT 4.400 94.840 496.000 96.240 ;
        RECT 4.000 88.080 496.000 94.840 ;
        RECT 4.400 86.680 496.000 88.080 ;
        RECT 4.000 79.920 496.000 86.680 ;
        RECT 4.400 78.520 496.000 79.920 ;
        RECT 4.000 71.760 496.000 78.520 ;
        RECT 4.400 70.360 496.000 71.760 ;
        RECT 4.000 68.360 496.000 70.360 ;
        RECT 4.000 66.960 495.600 68.360 ;
        RECT 4.000 62.920 496.000 66.960 ;
        RECT 4.400 61.520 496.000 62.920 ;
        RECT 4.000 54.760 496.000 61.520 ;
        RECT 4.400 53.360 496.000 54.760 ;
        RECT 4.000 46.600 496.000 53.360 ;
        RECT 4.400 45.200 496.000 46.600 ;
        RECT 4.000 38.440 496.000 45.200 ;
        RECT 4.400 37.040 496.000 38.440 ;
        RECT 4.000 29.600 496.000 37.040 ;
        RECT 4.400 28.200 496.000 29.600 ;
        RECT 4.000 23.480 496.000 28.200 ;
        RECT 4.000 22.080 495.600 23.480 ;
        RECT 4.000 21.440 496.000 22.080 ;
        RECT 4.400 20.040 496.000 21.440 ;
        RECT 4.000 13.280 496.000 20.040 ;
        RECT 4.400 11.880 496.000 13.280 ;
        RECT 4.000 5.120 496.000 11.880 ;
        RECT 4.400 4.255 496.000 5.120 ;
      LAYER met4 ;
        RECT 34.335 13.095 97.440 483.305 ;
        RECT 99.840 13.095 174.240 483.305 ;
        RECT 176.640 13.095 251.040 483.305 ;
        RECT 253.440 13.095 326.305 483.305 ;
  END
END Motor_Top
END LIBRARY

