* NGSPICE file created from Core.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

.subckt Core clock io_dbus_addr[0] io_dbus_addr[10] io_dbus_addr[11] io_dbus_addr[12]
+ io_dbus_addr[13] io_dbus_addr[14] io_dbus_addr[15] io_dbus_addr[16] io_dbus_addr[17]
+ io_dbus_addr[18] io_dbus_addr[19] io_dbus_addr[1] io_dbus_addr[20] io_dbus_addr[21]
+ io_dbus_addr[22] io_dbus_addr[23] io_dbus_addr[24] io_dbus_addr[25] io_dbus_addr[26]
+ io_dbus_addr[27] io_dbus_addr[28] io_dbus_addr[29] io_dbus_addr[2] io_dbus_addr[30]
+ io_dbus_addr[31] io_dbus_addr[3] io_dbus_addr[4] io_dbus_addr[5] io_dbus_addr[6]
+ io_dbus_addr[7] io_dbus_addr[8] io_dbus_addr[9] io_dbus_ld_type[0] io_dbus_ld_type[1]
+ io_dbus_ld_type[2] io_dbus_rd_en io_dbus_rdata[0] io_dbus_rdata[10] io_dbus_rdata[11]
+ io_dbus_rdata[12] io_dbus_rdata[13] io_dbus_rdata[14] io_dbus_rdata[15] io_dbus_rdata[16]
+ io_dbus_rdata[17] io_dbus_rdata[18] io_dbus_rdata[19] io_dbus_rdata[1] io_dbus_rdata[20]
+ io_dbus_rdata[21] io_dbus_rdata[22] io_dbus_rdata[23] io_dbus_rdata[24] io_dbus_rdata[25]
+ io_dbus_rdata[26] io_dbus_rdata[27] io_dbus_rdata[28] io_dbus_rdata[29] io_dbus_rdata[2]
+ io_dbus_rdata[30] io_dbus_rdata[31] io_dbus_rdata[3] io_dbus_rdata[4] io_dbus_rdata[5]
+ io_dbus_rdata[6] io_dbus_rdata[7] io_dbus_rdata[8] io_dbus_rdata[9] io_dbus_st_type[0]
+ io_dbus_st_type[1] io_dbus_valid io_dbus_wdata[0] io_dbus_wdata[10] io_dbus_wdata[11]
+ io_dbus_wdata[12] io_dbus_wdata[13] io_dbus_wdata[14] io_dbus_wdata[15] io_dbus_wdata[16]
+ io_dbus_wdata[17] io_dbus_wdata[18] io_dbus_wdata[19] io_dbus_wdata[1] io_dbus_wdata[20]
+ io_dbus_wdata[21] io_dbus_wdata[22] io_dbus_wdata[23] io_dbus_wdata[24] io_dbus_wdata[25]
+ io_dbus_wdata[26] io_dbus_wdata[27] io_dbus_wdata[28] io_dbus_wdata[29] io_dbus_wdata[2]
+ io_dbus_wdata[30] io_dbus_wdata[31] io_dbus_wdata[3] io_dbus_wdata[4] io_dbus_wdata[5]
+ io_dbus_wdata[6] io_dbus_wdata[7] io_dbus_wdata[8] io_dbus_wdata[9] io_dbus_wr_en
+ io_ibus_addr[0] io_ibus_addr[10] io_ibus_addr[11] io_ibus_addr[12] io_ibus_addr[13]
+ io_ibus_addr[14] io_ibus_addr[15] io_ibus_addr[16] io_ibus_addr[17] io_ibus_addr[18]
+ io_ibus_addr[19] io_ibus_addr[1] io_ibus_addr[20] io_ibus_addr[21] io_ibus_addr[22]
+ io_ibus_addr[23] io_ibus_addr[24] io_ibus_addr[25] io_ibus_addr[26] io_ibus_addr[27]
+ io_ibus_addr[28] io_ibus_addr[29] io_ibus_addr[2] io_ibus_addr[30] io_ibus_addr[31]
+ io_ibus_addr[3] io_ibus_addr[4] io_ibus_addr[5] io_ibus_addr[6] io_ibus_addr[7]
+ io_ibus_addr[8] io_ibus_addr[9] io_ibus_inst[0] io_ibus_inst[10] io_ibus_inst[11]
+ io_ibus_inst[12] io_ibus_inst[13] io_ibus_inst[14] io_ibus_inst[15] io_ibus_inst[16]
+ io_ibus_inst[17] io_ibus_inst[18] io_ibus_inst[19] io_ibus_inst[1] io_ibus_inst[20]
+ io_ibus_inst[21] io_ibus_inst[22] io_ibus_inst[23] io_ibus_inst[24] io_ibus_inst[25]
+ io_ibus_inst[26] io_ibus_inst[27] io_ibus_inst[28] io_ibus_inst[29] io_ibus_inst[2]
+ io_ibus_inst[30] io_ibus_inst[31] io_ibus_inst[3] io_ibus_inst[4] io_ibus_inst[5]
+ io_ibus_inst[6] io_ibus_inst[7] io_ibus_inst[8] io_ibus_inst[9] io_ibus_valid io_irq_m1_irq
+ io_irq_m2_irq io_irq_m3_irq io_irq_spi_irq io_irq_uart_irq reset vccd1 vssd1
XFILLER_100_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10213__S0 _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09671_ _09671_/A _09671_/B vssd1 vssd1 vccd1 vccd1 _09671_/Y sky130_fd_sc_hd__nor2_1
X_18869_ _19326_/CLK _18869_/D vssd1 vssd1 vccd1 vccd1 _18869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13615__A _13615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17521__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11135__A _11135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10841__A1 _10837_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14165__B _14168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09105_ _11376_/A _11376_/C _11495_/B _11285_/A vssd1 vssd1 vccd1 vccd1 _09119_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_148_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10185__S _10185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09259__B _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16661__A _16661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09974__S _10075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12346__B2 _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09938_ _09969_/A _09938_/B vssd1 vssd1 vccd1 vccd1 _09938_/X sky130_fd_sc_hd__or2_1
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10204__S0 _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09869_ _09869_/A vssd1 vssd1 vccd1 vccd1 _09869_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_46_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ _11901_/A _11901_/C _19737_/Q vssd1 vssd1 vccd1 vccd1 _11902_/A sky130_fd_sc_hd__a21oi_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15599__A1 _15497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12880_ _12883_/B _12883_/C _12869_/X vssd1 vssd1 vccd1 vccd1 _12880_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _11831_/A vssd1 vssd1 vccd1 vccd1 _11831_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14271__A1 _18451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17431__S _17435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _14572_/B vssd1 vssd1 vccd1 vccd1 _14550_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _18348_/Q _18342_/Q _11444_/X _11721_/A vssd1 vssd1 vccd1 vccd1 _11762_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13501_/A vssd1 vssd1 vccd1 vccd1 _18408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10713_ _10713_/A vssd1 vssd1 vccd1 vccd1 _10713_/X sky130_fd_sc_hd__buf_4
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14023__A1 _14126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _18511_/Q _19749_/Q _14487_/S vssd1 vssd1 vccd1 vccd1 _14482_/A sky130_fd_sc_hd__mux2_1
X_11693_ _18564_/Q _11371_/Y _12277_/B _11692_/X vssd1 vssd1 vccd1 vccd1 _11693_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16220_ _16042_/X _19085_/Q _16224_/S vssd1 vssd1 vccd1 vccd1 _16221_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13432_ _13428_/X _13429_/X _13431_/X _12629_/S _19791_/Q vssd1 vssd1 vccd1 vccd1
+ _13432_/X sky130_fd_sc_hd__o32a_1
XANTENNA__11699__B _13667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10644_ _19251_/Q _19022_/Q _18953_/Q _19347_/Q _10631_/X _10634_/X vssd1 vssd1 vccd1
+ vccd1 _10645_/B sky130_fd_sc_hd__mux4_1
XFILLER_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16151_ _16151_/A vssd1 vssd1 vccd1 vccd1 _19050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13363_ _18644_/Q _13363_/B vssd1 vssd1 vccd1 vccd1 _13363_/X sky130_fd_sc_hd__or2_1
X_10575_ _18826_/Q _19380_/Q _19542_/Q _18794_/Q _11088_/S _10368_/A vssd1 vssd1 vccd1
+ vccd1 _10575_/X sky130_fd_sc_hd__mux4_2
XFILLER_154_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15102_ _15116_/A vssd1 vssd1 vccd1 vccd1 _15102_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_23_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12314_ _19753_/Q vssd1 vssd1 vccd1 vccd1 _12315_/A sky130_fd_sc_hd__inv_2
X_16082_ _16082_/A vssd1 vssd1 vccd1 vccd1 _19028_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13294_ _13217_/X _13284_/Y _13293_/X _13229_/X _18633_/Q vssd1 vssd1 vccd1 vccd1
+ _13294_/X sky130_fd_sc_hd__a32o_4
XFILLER_108_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15033_ _16832_/A vssd1 vssd1 vccd1 vccd1 _15033_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15187__A _16689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12245_ _12246_/A _12267_/C vssd1 vssd1 vccd1 vccd1 _12245_/X sky130_fd_sc_hd__or2_1
XFILLER_47_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09185__A _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19841_ _19851_/CLK _19841_/D vssd1 vssd1 vccd1 vccd1 _19841_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_122_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10443__S0 _09673_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ _14203_/A _12176_/B vssd1 vssd1 vccd1 vccd1 _12181_/A sky130_fd_sc_hd__xor2_1
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold3_A hold3/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11127_ _18439_/Q vssd1 vssd1 vccd1 vccd1 _11127_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19772_ _19779_/CLK _19772_/D vssd1 vssd1 vccd1 vccd1 _19772_/Q sky130_fd_sc_hd__dfxtp_1
X_16984_ _16835_/X _19399_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16985_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16510__S _16514_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15935_ _14996_/X _18969_/Q _15935_/S vssd1 vssd1 vccd1 vccd1 _15936_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11848__B1 _19735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18723_ _19631_/CLK _18723_/D vssd1 vssd1 vccd1 vccd1 _18723_/Q sky130_fd_sc_hd__dfxtp_1
X_11058_ _09407_/A _11049_/X _11053_/X _11057_/X _10944_/A vssd1 vssd1 vccd1 vccd1
+ _11058_/X sky130_fd_sc_hd__a311o_1
XFILLER_37_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15039__B1 _14737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10009_ _10022_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _10009_/X sky130_fd_sc_hd__or2_1
XFILLER_3_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09910__C1 _09249_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18654_ _19568_/CLK _18654_/D vssd1 vssd1 vccd1 vccd1 _18654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15866_ _15009_/X _18938_/Q _15874_/S vssd1 vssd1 vccd1 vccd1 _15867_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10778__B _10778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13154__B _13154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14817_ _14366_/X _14827_/C _14816_/Y vssd1 vssd1 vccd1 vccd1 _14817_/Y sky130_fd_sc_hd__a21oi_1
X_17605_ _19660_/Q _16844_/A _17605_/S vssd1 vssd1 vccd1 vccd1 _17606_/A sky130_fd_sc_hd__mux2_1
X_18585_ _18585_/CLK _18585_/D vssd1 vssd1 vccd1 vccd1 _18585_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14965__S _14997_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15797_ _15797_/A vssd1 vssd1 vccd1 vccd1 _18907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16746__A _16845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17536_ _17592_/A vssd1 vssd1 vccd1 vccd1 _17605_/S sky130_fd_sc_hd__buf_8
XFILLER_83_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14748_ _14815_/A vssd1 vssd1 vccd1 vccd1 _14945_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_33_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17467_ _17467_/A vssd1 vssd1 vccd1 vccd1 _19597_/D sky130_fd_sc_hd__clkbuf_1
X_14679_ _14696_/A vssd1 vssd1 vccd1 vccd1 _14694_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__14014__A1 _11846_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16418_ _19173_/Q _15574_/X _16424_/S vssd1 vssd1 vccd1 vccd1 _16419_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19206_ _19723_/CLK _19206_/D vssd1 vssd1 vccd1 vccd1 _19206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17398_ _16752_/X _19567_/Q _17402_/S vssd1 vssd1 vccd1 vccd1 _17399_/A sky130_fd_sc_hd__mux2_1
X_19137_ _19838_/CLK _19137_/D vssd1 vssd1 vccd1 vccd1 _19137_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09977__C1 _09763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15796__S _15802_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16349_ _16125_/X _19143_/Q _16351_/S vssd1 vssd1 vccd1 vccd1 _16350_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19068_ _19838_/CLK _19068_/D vssd1 vssd1 vccd1 vccd1 _19068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15514__A1 _15513_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18019_ _19792_/Q vssd1 vssd1 vccd1 vccd1 _18023_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12514__A _13171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12233__B _13615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17516__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16420__S _16424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09723_ _09723_/A vssd1 vssd1 vccd1 vccd1 _09723_/X sky130_fd_sc_hd__buf_4
XANTENNA__10969__A _10969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09654_ _10379_/A _09654_/B vssd1 vssd1 vccd1 vccd1 _09654_/X sky130_fd_sc_hd__or2_1
XFILLER_94_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09585_ _18878_/Q _19336_/Q _10125_/A vssd1 vssd1 vccd1 vccd1 _09585_/X sky130_fd_sc_hd__mux2_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11067__A1 _10774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14176__A _14178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12016__A0 _12013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12408__B _12408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10027__C1 _09249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17487__A _17533_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10360_ _10566_/A vssd1 vssd1 vccd1 vccd1 _10477_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10291_ _18833_/Q _19387_/Q _19549_/Q _18801_/Q _09342_/A _09603_/A vssd1 vssd1 vccd1
+ vccd1 _10292_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12424__A _12424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12030_ _12030_/A _12030_/B _11969_/A _12008_/A vssd1 vssd1 vccd1 vccd1 _12131_/B
+ sky130_fd_sc_hd__or4bb_2
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09733__A _11185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13981_ _13978_/X _13984_/B _13979_/X _13980_/X vssd1 vssd1 vccd1 vccd1 _13981_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14492__A1 _19754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15720_ _15720_/A vssd1 vssd1 vccd1 vccd1 _18873_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12932_ _18288_/Q _12932_/B vssd1 vssd1 vccd1 vccd1 _12935_/B sky130_fd_sc_hd__nor2_1
XANTENNA__16769__A0 _16768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _15651_/A vssd1 vssd1 vccd1 vccd1 _18842_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12863_ _18268_/Q _12863_/B _12863_/C vssd1 vssd1 vccd1 vccd1 _12864_/C sky130_fd_sc_hd__and3_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14696_/A vssd1 vssd1 vccd1 vccd1 _14624_/A sky130_fd_sc_hd__clkbuf_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11058__A1 _09407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18370_ _19755_/CLK _18370_/D vssd1 vssd1 vccd1 vccd1 _18370_/Q sky130_fd_sc_hd__dfxtp_1
X_11814_ _19734_/Q vssd1 vssd1 vccd1 vccd1 _11849_/A sky130_fd_sc_hd__buf_4
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _15582_/A vssd1 vssd1 vccd1 vccd1 _18813_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _19858_/Q _19857_/Q vssd1 vssd1 vccd1 vccd1 _18214_/C sky130_fd_sc_hd__and2_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16285__B _17064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17321_ _17389_/S vssd1 vssd1 vccd1 vccd1 _17330_/S sky130_fd_sc_hd__buf_2
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14533_ _18563_/Q _14559_/B vssd1 vssd1 vccd1 vccd1 _14533_/X sky130_fd_sc_hd__or2_1
XFILLER_15_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11745_ _11745_/A _11745_/B vssd1 vssd1 vccd1 vccd1 _11747_/A sky130_fd_sc_hd__and2_2
XFILLER_15_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11503__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17252_ _19502_/Q _16645_/X _17258_/S vssd1 vssd1 vccd1 vccd1 _17253_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10900__S1 _10713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14464_ _14464_/A vssd1 vssd1 vccd1 vccd1 _18503_/D sky130_fd_sc_hd__clkbuf_1
X_11676_ _11676_/A vssd1 vssd1 vccd1 vccd1 _15263_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10018__C1 _09135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16203_ _16125_/X _19074_/Q _16205_/S vssd1 vssd1 vccd1 vccd1 _16204_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13415_ _13415_/A _18649_/Q vssd1 vssd1 vccd1 vccd1 _13415_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11222__B _12500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17183_ _17183_/A vssd1 vssd1 vccd1 vccd1 _19481_/D sky130_fd_sc_hd__clkbuf_1
X_10627_ _10875_/A _10627_/B vssd1 vssd1 vccd1 vccd1 _10627_/X sky130_fd_sc_hd__or2_1
XFILLER_139_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09423__A1 _09814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14395_ _18477_/Q _18509_/Q _14395_/S vssd1 vssd1 vccd1 vccd1 _14396_/A sky130_fd_sc_hd__mux2_1
X_16134_ _16844_/A vssd1 vssd1 vccd1 vccd1 _16134_/X sky130_fd_sc_hd__clkbuf_1
X_13346_ _13297_/X _13337_/Y _13345_/X _13306_/X _18641_/Q vssd1 vssd1 vccd1 vccd1
+ _13346_/X sky130_fd_sc_hd__a32o_4
XFILLER_6_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10558_ _18595_/Q _19284_/Q _10558_/S vssd1 vssd1 vccd1 vccd1 _10559_/B sky130_fd_sc_hd__mux2_1
XFILLER_170_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16065_ _16064_/X _19023_/Q _16065_/S vssd1 vssd1 vccd1 vccd1 _16066_/A sky130_fd_sc_hd__mux2_1
X_13277_ _19837_/Q _12736_/X _13276_/X vssd1 vssd1 vccd1 vccd1 _14859_/D sky130_fd_sc_hd__a21o_1
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10489_ _10485_/X _10487_/X _10488_/X _10392_/A _09529_/X vssd1 vssd1 vccd1 vccd1
+ _10494_/B sky130_fd_sc_hd__o221a_1
X_15016_ _15037_/C _15016_/B vssd1 vssd1 vccd1 vccd1 _15016_/X sky130_fd_sc_hd__or2_1
X_12228_ _12493_/C _12345_/A _12227_/X vssd1 vssd1 vccd1 vccd1 _14227_/A sky130_fd_sc_hd__o21ai_4
XFILLER_97_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19824_ _19866_/CLK _19824_/D vssd1 vssd1 vccd1 vccd1 _19824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16240__S _16246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12159_ _12160_/A _13598_/A vssd1 vssd1 vccd1 vccd1 _12161_/A sky130_fd_sc_hd__and2_1
XFILLER_97_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19755_ _19755_/CLK _19755_/D vssd1 vssd1 vccd1 vccd1 _19755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16967_ _16809_/X _19391_/Q _16975_/S vssd1 vssd1 vccd1 vccd1 _16968_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14483__A1 _12246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13165__A _15254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18706_ _19712_/CLK _18706_/D vssd1 vssd1 vccd1 vccd1 _18706_/Q sky130_fd_sc_hd__dfxtp_1
X_15918_ _14908_/X _18961_/Q _15924_/S vssd1 vssd1 vccd1 vccd1 _15919_/A sky130_fd_sc_hd__mux2_1
X_16898_ _19361_/Q _16712_/X _16902_/S vssd1 vssd1 vccd1 vccd1 _16899_/A sky130_fd_sc_hd__mux2_1
X_19686_ _19686_/CLK _19686_/D vssd1 vssd1 vccd1 vccd1 _19686_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15849_ _15849_/A vssd1 vssd1 vccd1 vccd1 _18930_/D sky130_fd_sc_hd__clkbuf_1
X_18637_ _19081_/CLK _18637_/D vssd1 vssd1 vccd1 vccd1 _18637_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14235__A1 _14232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17071__S _17075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09370_ _09370_/A _09370_/B vssd1 vssd1 vccd1 vccd1 _09370_/Y sky130_fd_sc_hd__nand2_1
X_18568_ _18585_/CLK _18568_/D vssd1 vssd1 vccd1 vccd1 _18568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17519_ _17519_/A vssd1 vssd1 vccd1 vccd1 _19621_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18499_ _19693_/CLK _18499_/D vssd1 vssd1 vccd1 vccd1 _18499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10029__A _10029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16150__S _16150_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10699__A _10724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14474__A1 _19746_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09706_ _18779_/Q _19008_/Q _18939_/Q _19237_/Q _09692_/A _09704_/A vssd1 vssd1 vccd1
+ vccd1 _09707_/B sky130_fd_sc_hd__mux4_1
XANTENNA__17770__A _18489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09637_ _19430_/Q _19206_/Q _19723_/Q _19174_/Q _11153_/A _09636_/X vssd1 vssd1 vccd1
+ vccd1 _09638_/B sky130_fd_sc_hd__mux4_1
XFILLER_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09699__S _10256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09568_ _09772_/A _09568_/B vssd1 vssd1 vccd1 vccd1 _09568_/X sky130_fd_sc_hd__or2_1
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09499_ _10581_/S vssd1 vssd1 vccd1 vccd1 _10401_/A sky130_fd_sc_hd__buf_4
XFILLER_168_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11530_ _11470_/A _13521_/B _11530_/C vssd1 vssd1 vccd1 vccd1 _11538_/B sky130_fd_sc_hd__and3b_1
XANTENNA__10894__S0 _10711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16923__A0 _16743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11461_ input72/X vssd1 vssd1 vccd1 vccd1 _14601_/A sky130_fd_sc_hd__clkinv_2
XFILLER_109_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13201__A2 _13197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16325__S _16329_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13200_ _18355_/Q _13246_/B vssd1 vssd1 vccd1 vccd1 _13200_/X sky130_fd_sc_hd__or2_1
X_10412_ _10412_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _10413_/B sky130_fd_sc_hd__nor2_1
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11392_ _11722_/C _11723_/A vssd1 vssd1 vccd1 vccd1 _11716_/A sky130_fd_sc_hd__and2b_2
X_14180_ _14312_/A _14180_/B vssd1 vssd1 vccd1 vccd1 _14180_/X sky130_fd_sc_hd__or2_1
XFILLER_109_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13131_ _19856_/Q _12604_/A _12584_/A _19824_/Q vssd1 vssd1 vccd1 vccd1 _13131_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10343_ _10327_/A _10342_/X _09317_/A vssd1 vssd1 vccd1 vccd1 _10343_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input55_A io_ibus_inst[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062_ _18331_/Q vssd1 vssd1 vccd1 vccd1 _13067_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10274_ _09277_/A _10264_/X _10273_/X _09284_/A _18442_/Q vssd1 vssd1 vccd1 vccd1
+ _10299_/A sky130_fd_sc_hd__a32o_4
XFILLER_97_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10949__S1 _09481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ _12013_/A _12013_/B vssd1 vssd1 vccd1 vccd1 _12013_/X sky130_fd_sc_hd__xor2_4
X_17870_ _17874_/A _17870_/B vssd1 vssd1 vccd1 vccd1 _17871_/A sky130_fd_sc_hd__or2_1
XFILLER_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16821_ _16821_/A vssd1 vssd1 vccd1 vccd1 _19330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_181_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19539_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__16995__S _17003_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14465__A1 _12067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16752_ _16752_/A vssd1 vssd1 vccd1 vccd1 _16752_/X sky130_fd_sc_hd__clkbuf_2
X_19540_ _19540_/CLK _19540_/D vssd1 vssd1 vccd1 vccd1 _19540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13964_ _13964_/A vssd1 vssd1 vccd1 vccd1 _13964_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09567__S1 _09144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15703_ _15703_/A vssd1 vssd1 vccd1 vccd1 _18865_/D sky130_fd_sc_hd__clkbuf_1
X_12915_ _12925_/C _12919_/C _12869_/X vssd1 vssd1 vccd1 vccd1 _12915_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19471_ _19472_/CLK _19471_/D vssd1 vssd1 vccd1 vccd1 _19471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16683_ _16683_/A vssd1 vssd1 vccd1 vccd1 _16683_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13895_ _14037_/A vssd1 vssd1 vccd1 vccd1 _14182_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15404__S _15406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18422_ _18506_/CLK _18422_/D vssd1 vssd1 vccd1 vccd1 _18422_/Q sky130_fd_sc_hd__dfxtp_1
X_15634_ _18835_/Q _15548_/X _15636_/S vssd1 vssd1 vccd1 vccd1 _15635_/A sky130_fd_sc_hd__mux2_1
X_12846_ _18264_/Q vssd1 vssd1 vccd1 vccd1 _12850_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13425__C1 _13401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _18357_/CLK _18353_/D vssd1 vssd1 vccd1 vccd1 _18353_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _18808_/Q _15564_/X _15568_/S vssd1 vssd1 vccd1 vccd1 _15566_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17167__A0 _18434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12777_ _12777_/A _12777_/B vssd1 vssd1 vccd1 vccd1 _12778_/B sky130_fd_sc_hd__or2_2
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09644__A1 _09171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _17304_/A vssd1 vssd1 vccd1 vccd1 _17313_/S sky130_fd_sc_hd__buf_4
XFILLER_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14516_ _11468_/B _18526_/Q _14516_/S vssd1 vssd1 vccd1 vccd1 _14517_/B sky130_fd_sc_hd__mux2_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18284_ _19759_/CLK _18284_/D vssd1 vssd1 vccd1 vccd1 _18284_/Q sky130_fd_sc_hd__dfxtp_1
X_11728_ _18353_/Q _11726_/Y _11888_/C vssd1 vssd1 vccd1 vccd1 _11728_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15496_ _15496_/A vssd1 vssd1 vccd1 vccd1 _18786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17235_ _18454_/Q _13399_/X _17235_/S vssd1 vssd1 vccd1 vccd1 _17235_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14447_ _14447_/A vssd1 vssd1 vccd1 vccd1 _18495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11659_ _19730_/Q _11788_/B vssd1 vssd1 vccd1 vccd1 _11684_/A sky130_fd_sc_hd__or2_1
XFILLER_31_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12400__A0 _11200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17166_ _17166_/A vssd1 vssd1 vccd1 vccd1 _19476_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10637__S0 _10631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09638__A _10309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14378_ _18471_/Q _18503_/Q _14381_/S vssd1 vssd1 vccd1 vccd1 _14379_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12951__A1 _18293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16117_ _16115_/X _19039_/Q _16129_/S vssd1 vssd1 vccd1 vccd1 _16118_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13329_ _13329_/A _13329_/B vssd1 vssd1 vccd1 vccd1 _14958_/B sky130_fd_sc_hd__or2_1
XANTENNA__17855__A _17895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17097_ _16790_/X _19449_/Q _17097_/S vssd1 vssd1 vccd1 vccd1 _17098_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_134_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _18623_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_115_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16048_ _16758_/A vssd1 vssd1 vccd1 vccd1 _16048_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15375__A _15397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19807_ _19810_/CLK _19807_/D vssd1 vssd1 vccd1 vccd1 _19807_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17642__A1 _17641_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_149_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19699_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10190__A1 _11178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17999_ _17999_/A vssd1 vssd1 vccd1 vccd1 _18027_/A sky130_fd_sc_hd__buf_2
XFILLER_38_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19738_ _19738_/CLK _19738_/D vssd1 vssd1 vccd1 vccd1 _19738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_145_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19669_ _19687_/CLK _19669_/D vssd1 vssd1 vccd1 vccd1 _19669_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__14208__A1 _12185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12219__A0 _14211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15314__S _15322_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13623__A _14216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09422_ _19660_/Q _19077_/Q _19114_/Q _18720_/Q _09367_/S _09364_/A vssd1 vssd1 vccd1
+ vccd1 _09422_/X sky130_fd_sc_hd__mux4_1
XANTENNA__14759__A2 _14703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09353_ _09353_/A vssd1 vssd1 vccd1 vccd1 _10651_/A sky130_fd_sc_hd__buf_2
XANTENNA__10485__A_N _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09284_ _09284_/A vssd1 vssd1 vccd1 vccd1 _09285_/A sky130_fd_sc_hd__buf_2
XANTENNA__10876__S0 _10614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17330__A0 _16758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09797__S1 _09763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10800__S0 _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10222__A _10447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10961_ _19504_/Q _19118_/Q _19568_/Q _18724_/Q _10959_/X _10960_/X vssd1 vssd1 vccd1
+ vccd1 _10962_/B sky130_fd_sc_hd__mux4_1
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15224__S _15233_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ _12766_/A vssd1 vssd1 vccd1 vccd1 _13426_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17005__A _17062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13680_ _13678_/X _13679_/X _13757_/S vssd1 vssd1 vccd1 vccd1 _13680_/X sky130_fd_sc_hd__mux2_1
X_10892_ _10899_/A _10889_/X _10891_/X vssd1 vssd1 vccd1 vccd1 _10892_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11108__S1 _10390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12631_ _18075_/A _12518_/X _12522_/X _13033_/A _12630_/X vssd1 vssd1 vccd1 vccd1
+ _12632_/B sky130_fd_sc_hd__a221o_2
XFILLER_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15350_ _15350_/A vssd1 vssd1 vccd1 vccd1 _18724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12562_ _18340_/Q _13042_/A vssd1 vssd1 vccd1 vccd1 _12562_/X sky130_fd_sc_hd__or2_1
XFILLER_157_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10867__S0 _10664_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14301_ _13943_/A _14296_/Y _14300_/Y vssd1 vssd1 vccd1 vccd1 _14301_/Y sky130_fd_sc_hd__a21oi_1
X_11513_ _11513_/A vssd1 vssd1 vccd1 vccd1 _14584_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15281_ _18694_/Q _15155_/X _15289_/S vssd1 vssd1 vccd1 vccd1 _15282_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16372__A1 _15506_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12493_ _12495_/A _12495_/B _12493_/C vssd1 vssd1 vccd1 vccd1 _12494_/A sky130_fd_sc_hd__and3_1
X_17020_ _17020_/A vssd1 vssd1 vccd1 vccd1 _19414_/D sky130_fd_sc_hd__clkbuf_1
X_14232_ _12244_/B _14102_/X _14231_/X vssd1 vssd1 vccd1 vccd1 _14232_/X sky130_fd_sc_hd__a21bo_1
XFILLER_172_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_51_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19589_/CLK sky130_fd_sc_hd__clkbuf_16
X_11444_ _18343_/Q _18338_/Q _18337_/Q _18344_/Q vssd1 vssd1 vccd1 vccd1 _11444_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_144_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11197__B1 _09430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15894__S _15902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14163_ _14163_/A _14319_/B vssd1 vssd1 vccd1 vccd1 _14163_/Y sky130_fd_sc_hd__nor2_1
X_11375_ _11375_/A _11375_/B vssd1 vssd1 vccd1 vccd1 _11639_/A sky130_fd_sc_hd__or2_1
XFILLER_164_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13114_ _18349_/Q _13109_/X _13113_/Y vssd1 vssd1 vccd1 vccd1 _18349_/D sky130_fd_sc_hd__o21a_1
X_10326_ _19418_/Q _19194_/Q _19711_/Q _19162_/Q _10125_/A _09723_/A vssd1 vssd1 vccd1
+ vccd1 _10327_/B sky130_fd_sc_hd__mux4_1
XFILLER_140_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18971_ _19591_/CLK _18971_/D vssd1 vssd1 vccd1 vccd1 _18971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14094_ _13806_/A _14092_/B _14093_/X _14037_/A vssd1 vssd1 vccd1 vccd1 _14094_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15883__A0 _14714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_66_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19822_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _19821_/Q _19820_/Q _19822_/Q _18097_/A vssd1 vssd1 vccd1 vccd1 _17927_/D
+ sky130_fd_sc_hd__and4_1
X_13045_ _18326_/Q _13045_/B _13045_/C vssd1 vssd1 vccd1 vccd1 _13046_/C sky130_fd_sc_hd__and3_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10257_ _18865_/Q _19323_/Q _10257_/S vssd1 vssd1 vccd1 vccd1 _10257_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17624__A1 _17623_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10188_ _18771_/Q _19000_/Q _18931_/Q _19229_/Q _09721_/X _09723_/X vssd1 vssd1 vccd1
+ vccd1 _10188_/X sky130_fd_sc_hd__mux4_1
X_17853_ _15238_/X _19727_/Q _17853_/S vssd1 vssd1 vccd1 vccd1 _17854_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16804_ _16803_/X _19325_/Q _16807_/S vssd1 vssd1 vccd1 vccd1 _16805_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10132__A _10132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14996_ _16822_/A vssd1 vssd1 vccd1 vccd1 _14996_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17784_ _17840_/A vssd1 vssd1 vccd1 vccd1 _17853_/S sky130_fd_sc_hd__buf_6
XFILLER_82_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19523_ _19838_/CLK _19523_/D vssd1 vssd1 vccd1 vccd1 _19523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13947_ _14135_/A _13946_/Y _13816_/X vssd1 vssd1 vccd1 vccd1 _13947_/X sky130_fd_sc_hd__o21a_1
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16735_ _19304_/Q _16734_/X _16735_/S vssd1 vssd1 vccd1 vccd1 _16736_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11121__B1 _10219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19454_ _19584_/CLK _19454_/D vssd1 vssd1 vccd1 vccd1 _19454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16666_ _16666_/A vssd1 vssd1 vccd1 vccd1 _19282_/D sky130_fd_sc_hd__clkbuf_1
X_13878_ _13876_/X _13877_/X _13913_/S vssd1 vssd1 vccd1 vccd1 _13878_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18405_ _19689_/CLK _18405_/D vssd1 vssd1 vccd1 vccd1 _18405_/Q sky130_fd_sc_hd__dfxtp_1
X_15617_ _18827_/Q _15522_/X _15625_/S vssd1 vssd1 vccd1 vccd1 _15618_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12829_ _12830_/B _12830_/C _18259_/Q vssd1 vssd1 vccd1 vccd1 _12831_/B sky130_fd_sc_hd__a21oi_1
X_16597_ _19254_/Q vssd1 vssd1 vccd1 vccd1 _16598_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_50_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19385_ _19579_/CLK _19385_/D vssd1 vssd1 vccd1 vccd1 _19385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09617__A1 _11178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18336_ _18401_/CLK _18336_/D vssd1 vssd1 vccd1 vccd1 _18336_/Q sky130_fd_sc_hd__dfxtp_1
X_15548_ _16803_/A vssd1 vssd1 vccd1 vccd1 _15548_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18267_ _19779_/CLK _18267_/D vssd1 vssd1 vccd1 vccd1 _18267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15479_ _18781_/Q _15229_/X _15481_/S vssd1 vssd1 vccd1 vccd1 _15480_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16363__A1 _15494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14274__A _14274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_19_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19713_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_163_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17218_ _18449_/Q _12757_/X _17218_/S vssd1 vssd1 vccd1 vccd1 _17218_/X sky130_fd_sc_hd__mux2_1
X_18198_ _19853_/Q _18194_/B _18197_/Y vssd1 vssd1 vccd1 vccd1 _19853_/D sky130_fd_sc_hd__o21a_1
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_71_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17149_ _17762_/S _17149_/B vssd1 vssd1 vccd1 vccd1 _17149_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09250__C1 _09249_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09971_ _09879_/A _09970_/X _09319_/A vssd1 vssd1 vccd1 vccd1 _09971_/X sky130_fd_sc_hd__o21a_1
XFILLER_118_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15309__S _15311_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12522__A _12602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14168__B _14168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09405_ _18980_/Q vssd1 vssd1 vccd1 vccd1 _10774_/A sky130_fd_sc_hd__inv_2
XFILLER_38_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15979__S _15983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16664__A _16664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09336_ _09336_/A vssd1 vssd1 vccd1 vccd1 _10706_/S sky130_fd_sc_hd__buf_6
XANTENNA__10849__S0 _10648_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09267_ _16212_/A _18570_/Q vssd1 vssd1 vccd1 vccd1 _09267_/X sky130_fd_sc_hd__or2b_1
XANTENNA__13168__A1 _13139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09198_ _11097_/A vssd1 vssd1 vccd1 vccd1 _09640_/A sky130_fd_sc_hd__buf_2
XFILLER_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09241__C1 _09231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11160_ _19431_/Q _19207_/Q _19724_/Q _19175_/Q _11153_/X _09542_/A vssd1 vssd1 vccd1
+ vccd1 _11160_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14668__A1 _14568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14668__B2 input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10111_ _10107_/A _10108_/X _10110_/X _09988_/X vssd1 vssd1 vccd1 vccd1 _10111_/X
+ sky130_fd_sc_hd__o211a_1
X_11091_ _19416_/Q _19192_/Q _19709_/Q _19160_/Q _10348_/S _09539_/A vssd1 vssd1 vccd1
+ vccd1 _11091_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12432__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10042_ _10042_/A _10042_/B vssd1 vssd1 vccd1 vccd1 _10042_/X sky130_fd_sc_hd__or2_1
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13962__S _14032_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14850_ _18438_/Q _12726_/B _15051_/S vssd1 vssd1 vccd1 vccd1 _14850_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13801_ _13801_/A vssd1 vssd1 vccd1 vccd1 _14040_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14781_ _16661_/A vssd1 vssd1 vccd1 vccd1 _16765_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input18_A io_dbus_rdata[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ _13265_/A _12020_/C vssd1 vssd1 vccd1 vccd1 _11993_/X sky130_fd_sc_hd__or2_1
XANTENNA__10887__A _10887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16520_ _16520_/A vssd1 vssd1 vccd1 vccd1 _19217_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13732_ _13922_/A _13729_/B vssd1 vssd1 vccd1 vccd1 _13870_/A sky130_fd_sc_hd__or2b_1
X_10944_ _10944_/A _10944_/B _10944_/C vssd1 vssd1 vccd1 vccd1 _10944_/X sky130_fd_sc_hd__or3_1
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15889__S _15891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16451_ _16061_/X _19187_/Q _16453_/S vssd1 vssd1 vccd1 vccd1 _16452_/A sky130_fd_sc_hd__mux2_1
X_13663_ _13661_/X _13662_/X _13742_/S vssd1 vssd1 vccd1 vccd1 _13663_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10875_ _10875_/A _10875_/B vssd1 vssd1 vccd1 vccd1 _10875_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14793__S _14822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15402_ _18748_/Q _15226_/X _15406_/S vssd1 vssd1 vccd1 vccd1 _15403_/A sky130_fd_sc_hd__mux2_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19170_ _19557_/CLK _19170_/D vssd1 vssd1 vccd1 vccd1 _19170_/Q sky130_fd_sc_hd__dfxtp_1
X_12614_ _19810_/Q _12518_/A _12602_/X _18321_/Q _12613_/X vssd1 vssd1 vccd1 vccd1
+ _12615_/B sky130_fd_sc_hd__a221o_2
X_16382_ _16428_/S vssd1 vssd1 vccd1 vccd1 _16391_/S sky130_fd_sc_hd__buf_2
X_13594_ _13594_/A vssd1 vssd1 vccd1 vccd1 _13594_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18121_ _18199_/A vssd1 vssd1 vccd1 vccd1 _18159_/A sky130_fd_sc_hd__clkbuf_2
X_15333_ _18718_/Q _15232_/X _15333_/S vssd1 vssd1 vccd1 vccd1 _15334_/A sky130_fd_sc_hd__mux2_1
X_12545_ _12545_/A _12567_/A vssd1 vssd1 vccd1 vccd1 _12546_/A sky130_fd_sc_hd__and2_1
XFILLER_12_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18052_ _18051_/B _18051_/C _19803_/Q vssd1 vssd1 vccd1 vccd1 _18053_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__11511__A _11511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15264_ _18688_/Q _15263_/X _15264_/S vssd1 vssd1 vccd1 vccd1 _15265_/A sky130_fd_sc_hd__mux2_1
X_12476_ _12472_/A _12476_/B vssd1 vssd1 vccd1 vccd1 _12477_/A sky130_fd_sc_hd__and2b_1
XFILLER_144_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17003_ _19407_/Q _16654_/X _17003_/S vssd1 vssd1 vccd1 vccd1 _17004_/A sky130_fd_sc_hd__mux2_1
X_14215_ _14323_/A _14215_/B vssd1 vssd1 vccd1 vccd1 _14215_/Y sky130_fd_sc_hd__nor2_1
X_11427_ _11427_/A _11427_/B _12516_/A _15241_/A vssd1 vssd1 vccd1 vccd1 _11427_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__09232__C1 _09231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ _18668_/Q _15194_/X _15201_/S vssd1 vssd1 vccd1 vccd1 _15196_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14146_ _13949_/A _14143_/X _14145_/Y _13726_/X vssd1 vssd1 vccd1 vccd1 _14146_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_152_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11358_ _11361_/A _11358_/B _11642_/C vssd1 vssd1 vccd1 vccd1 _11584_/A sky130_fd_sc_hd__nor3_2
XFILLER_98_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10881__A2_N _10834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10309_ _10309_/A _10309_/B vssd1 vssd1 vccd1 vccd1 _10309_/X sky130_fd_sc_hd__or2_1
X_18954_ _19726_/CLK _18954_/D vssd1 vssd1 vccd1 vccd1 _18954_/Q sky130_fd_sc_hd__dfxtp_1
X_14077_ _13927_/A _14078_/B _14076_/X _13856_/A vssd1 vssd1 vccd1 vccd1 _14077_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_98_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11289_ _11279_/Y _11281_/Y _11284_/Y _11286_/X _11288_/X vssd1 vssd1 vccd1 vccd1
+ _11565_/B sky130_fd_sc_hd__o2111a_1
X_17905_ _19754_/Q _17886_/X _12339_/X _12342_/Y _17895_/X vssd1 vssd1 vccd1 vccd1
+ _19754_/D sky130_fd_sc_hd__o221a_1
X_13028_ _13049_/A _13033_/C vssd1 vssd1 vccd1 vccd1 _13028_/Y sky130_fd_sc_hd__nor2_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18885_ _19700_/CLK _18885_/D vssd1 vssd1 vccd1 vccd1 _18885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17344__S _17352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17836_ _15213_/X _19719_/Q _17838_/S vssd1 vssd1 vccd1 vccd1 _17837_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09651__A _10309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17767_ _17770_/B _17766_/Y _17713_/X vssd1 vssd1 vccd1 vccd1 _17767_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10797__A _10797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14979_ _18480_/Q _18481_/Q _14979_/C vssd1 vssd1 vccd1 vccd1 _15002_/C sky130_fd_sc_hd__and3_1
X_19506_ _19506_/CLK _19506_/D vssd1 vssd1 vccd1 vccd1 _19506_/Q sky130_fd_sc_hd__dfxtp_1
X_16718_ _16718_/A vssd1 vssd1 vccd1 vccd1 _16718_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17698_ _12598_/B _17697_/Y _17734_/S vssd1 vssd1 vccd1 vccd1 _17698_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11197__A1_N _18454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19437_ _19599_/CLK _19437_/D vssd1 vssd1 vccd1 vccd1 _19437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16649_ _19277_/Q _16648_/X _16655_/S vssd1 vssd1 vccd1 vccd1 _16650_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19368_ _19626_/CLK _19368_/D vssd1 vssd1 vccd1 vccd1 _19368_/Q sky130_fd_sc_hd__dfxtp_1
X_09121_ _18555_/Q vssd1 vssd1 vccd1 vccd1 _11297_/B sky130_fd_sc_hd__clkbuf_1
X_18319_ _19812_/CLK _18319_/D vssd1 vssd1 vccd1 vccd1 _18319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19299_ _19395_/CLK _19299_/D vssd1 vssd1 vccd1 vccd1 _19299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14732__A _14842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09826__A _09826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12373__A2 _14289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11581__B1 _18574_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09954_ _19329_/Q vssd1 vssd1 vccd1 vccd1 _09954_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09885_ _19622_/Q _19460_/Q _18906_/Q _18676_/Q _09866_/X _09869_/X vssd1 vssd1 vccd1
+ vccd1 _09886_/B sky130_fd_sc_hd__mux4_1
XFILLER_100_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17254__S _17258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11636__A1 _14555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10500__A _10500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11100__A3 _18798_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17772__A0 _19690_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14907__A _16693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10660_ _11077_/A _12473_/A vssd1 vssd1 vccd1 vccd1 _11080_/B sky130_fd_sc_hd__nand2_1
XFILLER_41_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09500__S _10401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09319_ _09319_/A vssd1 vssd1 vccd1 vccd1 _09320_/A sky130_fd_sc_hd__buf_2
X_10591_ _10591_/A _10591_/B vssd1 vssd1 vccd1 vccd1 _10591_/X sky130_fd_sc_hd__or2_1
XFILLER_167_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10072__B1 _09309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12330_ _12330_/A _12355_/A vssd1 vssd1 vccd1 vccd1 _12371_/B sky130_fd_sc_hd__xor2_4
XFILLER_126_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11688__D _13845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17429__S _17435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15738__A _15806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ _12286_/A vssd1 vssd1 vccd1 vccd1 _12262_/B sky130_fd_sc_hd__clkinv_4
XFILLER_135_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14000_ _14037_/A vssd1 vssd1 vccd1 vccd1 _14000_/X sky130_fd_sc_hd__clkbuf_2
X_11212_ _11321_/C _14519_/A _11534_/B vssd1 vssd1 vccd1 vccd1 _11299_/A sky130_fd_sc_hd__nand3b_1
XFILLER_134_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12192_ _19679_/Q _13529_/B vssd1 vssd1 vccd1 vccd1 _12192_/X sky130_fd_sc_hd__or2_1
XFILLER_123_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13258__A _18629_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11143_ _11227_/A _11229_/A _11227_/C _10102_/A _11142_/Y vssd1 vssd1 vccd1 vccd1
+ _11269_/C sky130_fd_sc_hd__a311o_1
XFILLER_150_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput75 _11956_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[11] sky130_fd_sc_hd__buf_2
XANTENNA__13313__A1 _12559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput86 _12213_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[21] sky130_fd_sc_hd__buf_2
Xoutput97 _12450_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[31] sky130_fd_sc_hd__buf_2
X_15951_ _15951_/A vssd1 vssd1 vccd1 vccd1 _18976_/D sky130_fd_sc_hd__clkbuf_1
X_11074_ _10691_/X _12469_/A _11779_/A _12466_/A vssd1 vssd1 vccd1 vccd1 _11257_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10025_ _10074_/A _10025_/B vssd1 vssd1 vccd1 vccd1 _10025_/X sky130_fd_sc_hd__or2_1
X_14902_ _14802_/A _14802_/B _11305_/A input7/X _14803_/B vssd1 vssd1 vccd1 vccd1
+ _15000_/A sky130_fd_sc_hd__a41o_1
X_18670_ _19165_/CLK _18670_/D vssd1 vssd1 vccd1 vccd1 _18670_/Q sky130_fd_sc_hd__dfxtp_1
X_15882_ _15950_/S vssd1 vssd1 vccd1 vccd1 _15891_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_48_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11875__B2 _13658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17621_ _17621_/A _18462_/Q _17621_/C vssd1 vssd1 vccd1 vccd1 _17632_/C sky130_fd_sc_hd__or3_4
X_14833_ _16777_/A vssd1 vssd1 vccd1 vccd1 _14833_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14089__A _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17552_ _17552_/A vssd1 vssd1 vccd1 vccd1 _19635_/D sky130_fd_sc_hd__clkbuf_1
X_14764_ _14765_/A _14765_/C _17632_/A vssd1 vssd1 vccd1 vccd1 _14766_/A sky130_fd_sc_hd__a21oi_1
X_11976_ _11919_/A _11952_/A _11954_/B vssd1 vssd1 vccd1 vccd1 _11976_/Y sky130_fd_sc_hd__a21oi_1
X_16503_ _16503_/A _16503_/B vssd1 vssd1 vccd1 vccd1 _16560_/A sky130_fd_sc_hd__nor2_2
X_13715_ _14274_/A vssd1 vssd1 vccd1 vccd1 _14332_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10927_ _19599_/Q _19437_/Q _18883_/Q _18653_/Q _10959_/A _10960_/A vssd1 vssd1 vccd1
+ vccd1 _10928_/B sky130_fd_sc_hd__mux4_1
X_17483_ _19605_/Q _16667_/X _17485_/S vssd1 vssd1 vccd1 vccd1 _17484_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17763__A0 _19688_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14695_ _14695_/A vssd1 vssd1 vccd1 vccd1 _18584_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16508__S _16514_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19222_ _19707_/CLK _19222_/D vssd1 vssd1 vccd1 vccd1 _19222_/Q sky130_fd_sc_hd__dfxtp_1
X_13646_ _13667_/A _12381_/A _13659_/S vssd1 vssd1 vccd1 vccd1 _13646_/X sky130_fd_sc_hd__mux2_1
X_16434_ _16033_/X _19179_/Q _16442_/S vssd1 vssd1 vccd1 vccd1 _16435_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10858_ _10858_/A _18854_/Q vssd1 vssd1 vccd1 vccd1 _10858_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _19149_/Q _15497_/X _16369_/S vssd1 vssd1 vccd1 vccd1 _16366_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19153_ _19702_/CLK _19153_/D vssd1 vssd1 vccd1 vccd1 _19153_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10289__S1 _10239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13577_ _11551_/A _11333_/X _11476_/B _11531_/X _13520_/A vssd1 vssd1 vccd1 vccd1
+ _13579_/C sky130_fd_sc_hd__o311ai_1
X_10789_ _18853_/Q _19311_/Q _10886_/S vssd1 vssd1 vccd1 vccd1 _10790_/B sky130_fd_sc_hd__mux2_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18104_ _18120_/A _18104_/B _18104_/C vssd1 vssd1 vccd1 vccd1 _19821_/D sky130_fd_sc_hd__nor3_1
X_15316_ _18710_/Q _15207_/X _15322_/S vssd1 vssd1 vccd1 vccd1 _15317_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14329__B1 _15123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12528_ _12528_/A vssd1 vssd1 vccd1 vccd1 _12528_/X sky130_fd_sc_hd__clkbuf_2
X_16296_ _16048_/X _19119_/Q _16296_/S vssd1 vssd1 vccd1 vccd1 _16297_/A sky130_fd_sc_hd__mux2_1
X_19084_ _19630_/CLK _19084_/D vssd1 vssd1 vccd1 vccd1 _19084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15247_ _15247_/A vssd1 vssd1 vccd1 vccd1 _18683_/D sky130_fd_sc_hd__clkbuf_1
X_18035_ _18199_/A vssd1 vssd1 vccd1 vccd1 _18071_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12459_ _12459_/A vssd1 vssd1 vccd1 vccd1 _12459_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15178_ _16680_/A vssd1 vssd1 vccd1 vccd1 _15178_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09851__S0 _10010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14129_ _14124_/A _14126_/B _13795_/A _14127_/X _14128_/X vssd1 vssd1 vccd1 vccd1
+ _14130_/B sky130_fd_sc_hd__o221a_1
XFILLER_99_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18937_ _19557_/CLK _18937_/D vssd1 vssd1 vccd1 vccd1 _18937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10213__S1 _10080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _19270_/Q _19041_/Q _18972_/Q _19366_/Q _09600_/A _09603_/A vssd1 vssd1 vccd1
+ vccd1 _09671_/B sky130_fd_sc_hd__mux4_1
X_18868_ _19553_/CLK _18868_/D vssd1 vssd1 vccd1 vccd1 _18868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17819_ _15187_/X _19711_/Q _17827_/S vssd1 vssd1 vccd1 vccd1 _17820_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18799_ _19223_/CLK _18799_/D vssd1 vssd1 vccd1 vccd1 _18799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09906__S1 _09783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10320__A _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11135__B _12483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16418__S _16424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15322__S _15322_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_15_0_clock clkbuf_3_7_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_15_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10466__S _10466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09104_ _11317_/A _11325_/C vssd1 vssd1 vccd1 vccd1 _11285_/A sky130_fd_sc_hd__and2_1
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09937_ _18776_/Q _19005_/Q _18936_/Q _19234_/Q _09803_/A _09936_/X vssd1 vssd1 vccd1
+ vccd1 _09938_/B sky130_fd_sc_hd__mux4_1
XFILLER_77_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09868_ _10029_/A vssd1 vssd1 vccd1 vccd1 _09869_/A sky130_fd_sc_hd__buf_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10204__S1 _10080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13525__B _14431_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _09788_/A _09791_/X _09798_/X _09231_/A vssd1 vssd1 vccd1 vccd1 _09799_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_46_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11830_ _11849_/A _11705_/X _11819_/X _11829_/X vssd1 vssd1 vccd1 vccd1 _17866_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13244__C _14813_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _18415_/Q _11022_/X _11716_/A _11676_/A vssd1 vssd1 vccd1 vccd1 _11764_/A
+ sky130_fd_sc_hd__a211o_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _18408_/Q _13364_/X _13508_/S vssd1 vssd1 vccd1 vccd1 _13501_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _10712_/A vssd1 vssd1 vccd1 vccd1 _10713_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14480_/A vssd1 vssd1 vccd1 vccd1 _18510_/D sky130_fd_sc_hd__clkbuf_1
X_11692_ _11692_/A _11692_/B _11692_/C vssd1 vssd1 vccd1 vccd1 _11692_/X sky130_fd_sc_hd__or3_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13431_ _18298_/Q _13404_/B _12703_/A _19690_/Q _13430_/X vssd1 vssd1 vccd1 vccd1
+ _13431_/X sky130_fd_sc_hd__a221o_1
X_10643_ _09409_/A _10636_/Y _10638_/Y _10640_/Y _10642_/Y vssd1 vssd1 vccd1 vccd1
+ _10643_/X sky130_fd_sc_hd__o32a_1
XFILLER_167_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12157__A _14192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16150_ _16048_/X _19050_/Q _16150_/S vssd1 vssd1 vccd1 vccd1 _16151_/A sky130_fd_sc_hd__mux2_1
X_13362_ _19785_/Q _13123_/X _13358_/X _13361_/X vssd1 vssd1 vccd1 vccd1 _13363_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_139_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10574_ _10574_/A _10574_/B vssd1 vssd1 vccd1 vccd1 _10574_/X sky130_fd_sc_hd__or2_1
XFILLER_166_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15101_ _18627_/Q _13566_/X _15097_/X _11077_/A vssd1 vssd1 vccd1 vccd1 _18627_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12313_ _12313_/A _12313_/B vssd1 vssd1 vccd1 vccd1 _12313_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__12591__S _12628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16081_ _16080_/X _19028_/Q _16081_/S vssd1 vssd1 vccd1 vccd1 _16082_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13293_ _18633_/Q _14873_/B _14873_/C _14873_/D vssd1 vssd1 vccd1 vccd1 _13293_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15032_ _16728_/A vssd1 vssd1 vccd1 vccd1 _16832_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12244_ _12411_/B _12244_/B vssd1 vssd1 vccd1 vccd1 _12244_/X sky130_fd_sc_hd__and2b_1
XFILLER_135_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14091__B _14093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19840_ _19851_/CLK _19840_/D vssd1 vssd1 vccd1 vccd1 _19840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10443__S1 _09486_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12175_ _12129_/A _12132_/B _14192_/A _12057_/A vssd1 vssd1 vccd1 vccd1 _12176_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_123_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15287__A1 _15165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11126_ _11119_/Y _11121_/Y _11123_/Y _11125_/Y _10494_/A vssd1 vssd1 vccd1 vccd1
+ _11126_/X sky130_fd_sc_hd__o221a_2
X_19771_ _19779_/CLK _19771_/D vssd1 vssd1 vccd1 vccd1 _19771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16983_ _16983_/A vssd1 vssd1 vccd1 vccd1 _19398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18722_ _19630_/CLK _18722_/D vssd1 vssd1 vccd1 vccd1 _18722_/Q sky130_fd_sc_hd__dfxtp_1
X_15934_ _15934_/A vssd1 vssd1 vccd1 vccd1 _18968_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11848__A1 _11849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ _10797_/A _11054_/X _11056_/X _10728_/A vssd1 vssd1 vccd1 vccd1 _11057_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10008_ _19264_/Q _19035_/Q _18966_/Q _19360_/Q _10075_/S _09147_/A vssd1 vssd1 vccd1
+ vccd1 _10009_/B sky130_fd_sc_hd__mux4_1
XFILLER_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13435__B _13435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18653_ _19698_/CLK _18653_/D vssd1 vssd1 vccd1 vccd1 _18653_/Q sky130_fd_sc_hd__dfxtp_1
X_15865_ _15865_/A vssd1 vssd1 vccd1 vccd1 _15874_/S sky130_fd_sc_hd__buf_4
XFILLER_36_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14798__A0 _18434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17604_ _17604_/A vssd1 vssd1 vccd1 vccd1 _19659_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14816_ _14366_/X _14827_/C _14829_/B vssd1 vssd1 vccd1 vccd1 _14816_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_36_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18584_ _18585_/CLK _18584_/D vssd1 vssd1 vccd1 vccd1 _18584_/Q sky130_fd_sc_hd__dfxtp_1
X_15796_ _15022_/X _18907_/Q _15802_/S vssd1 vssd1 vccd1 vccd1 _15797_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17535_ _17535_/A _17535_/B vssd1 vssd1 vccd1 vccd1 _17592_/A sky130_fd_sc_hd__nor2_4
XFILLER_45_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11959_ _19670_/Q _11959_/B vssd1 vssd1 vccd1 vccd1 _11959_/X sky130_fd_sc_hd__or2_1
XFILLER_17_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14747_ _18429_/Q _15071_/S vssd1 vssd1 vccd1 vccd1 _14747_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__16238__S _16246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10284__B1 _09315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17466_ _19597_/Q _16639_/X _17474_/S vssd1 vssd1 vccd1 vccd1 _17467_/A sky130_fd_sc_hd__mux2_1
X_14678_ _14678_/A vssd1 vssd1 vccd1 vccd1 _18579_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19205_ _19722_/CLK _19205_/D vssd1 vssd1 vccd1 vccd1 _19205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13222__A0 _11406_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16417_ _16417_/A vssd1 vssd1 vccd1 vccd1 _19172_/D sky130_fd_sc_hd__clkbuf_1
X_13629_ _13613_/X _13627_/X _13991_/S vssd1 vssd1 vccd1 vccd1 _13629_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17397_ _17397_/A vssd1 vssd1 vccd1 vccd1 _19566_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16762__A _16845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19136_ _19818_/CLK _19136_/D vssd1 vssd1 vccd1 vccd1 _19136_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14970__A0 _18448_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16348_ _16348_/A vssd1 vssd1 vccd1 vccd1 _19142_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17069__S _17075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19067_ _19812_/CLK _19067_/D vssd1 vssd1 vccd1 vccd1 _19067_/Q sky130_fd_sc_hd__dfxtp_1
X_16279_ _16128_/X _19112_/Q _16279_/S vssd1 vssd1 vccd1 vccd1 _16280_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10682__S1 _09139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18018_ _19791_/Q _18015_/B _18017_/Y vssd1 vssd1 vccd1 vccd1 _19791_/D sky130_fd_sc_hd__o21a_1
XANTENNA__09376__A _10950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09722_ _10280_/A vssd1 vssd1 vccd1 vccd1 _09723_/A sky130_fd_sc_hd__buf_2
XFILLER_101_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10198__S0 _10094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13345__B _13345_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ _18844_/Q _19398_/Q _19560_/Q _18812_/Q _09448_/S _10349_/A vssd1 vssd1 vccd1
+ vccd1 _09654_/B sky130_fd_sc_hd__mux4_1
XFILLER_95_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09584_ _10328_/S vssd1 vssd1 vccd1 vccd1 _10125_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16148__S _16150_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10370__S0 _09631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14176__B _14176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14891__S _14941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10578__B2 _18435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14192__A _14192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10290_ _11123_/A _10289_/X _09412_/A vssd1 vssd1 vccd1 vccd1 _10290_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09815__S0 _09803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15227__S _15233_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13536__A _13536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13980_ _14332_/A _13984_/A vssd1 vssd1 vccd1 vccd1 _13980_/X sky130_fd_sc_hd__or2_1
XFILLER_101_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10189__S0 _10129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12931_ _12943_/A _12931_/B _12932_/B vssd1 vssd1 vccd1 vccd1 _18287_/D sky130_fd_sc_hd__nor3_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16847__A _16847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17442__S _17446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12862_ _12863_/B _12863_/C _18268_/Q vssd1 vssd1 vccd1 vccd1 _12864_/B sky130_fd_sc_hd__a21oi_1
XFILLER_160_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _18842_/Q _15570_/X _15658_/S vssd1 vssd1 vccd1 vccd1 _15651_/A sky130_fd_sc_hd__mux2_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _14601_/A vssd1 vssd1 vccd1 vccd1 _14696_/A sky130_fd_sc_hd__clkbuf_2
X_11813_ _11844_/B _11813_/B vssd1 vssd1 vccd1 vccd1 _11813_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_33_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _18813_/Q _15580_/X _15584_/S vssd1 vssd1 vccd1 vccd1 _15582_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17718__A0 _19679_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12255__A1 _12495_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12793_ _11462_/A _13532_/A _18205_/B _19856_/Q vssd1 vssd1 vccd1 vccd1 _18214_/B
+ sky130_fd_sc_hd__and4bb_4
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09656__C1 _09247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _17376_/A vssd1 vssd1 vccd1 vccd1 _17389_/S sky130_fd_sc_hd__buf_8
X_14532_ _14565_/A vssd1 vssd1 vccd1 vccd1 _14559_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _11785_/A _11784_/A vssd1 vssd1 vccd1 vccd1 _11745_/B sky130_fd_sc_hd__or2_1
XFILLER_18_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17251_ _17251_/A vssd1 vssd1 vccd1 vccd1 _19501_/D sky130_fd_sc_hd__clkbuf_1
X_14463_ _18503_/Q _12043_/A _14465_/S vssd1 vssd1 vccd1 vccd1 _14464_/A sky130_fd_sc_hd__mux2_1
X_11675_ _11672_/Y _11674_/X _11720_/A vssd1 vssd1 vccd1 vccd1 _11678_/B sky130_fd_sc_hd__a21oi_2
XFILLER_168_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13414_ _13354_/X _13412_/X _13413_/X _13401_/X vssd1 vssd1 vccd1 vccd1 _18379_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09895__S _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16202_ _16202_/A vssd1 vssd1 vccd1 vccd1 _19073_/D sky130_fd_sc_hd__clkbuf_1
X_17182_ _19481_/Q _17181_/X _17189_/S vssd1 vssd1 vccd1 vccd1 _17183_/A sky130_fd_sc_hd__mux2_1
X_10626_ _19605_/Q _19443_/Q _18889_/Q _18659_/Q _10733_/S _10548_/A vssd1 vssd1 vccd1
+ vccd1 _10627_/B sky130_fd_sc_hd__mux4_1
XFILLER_167_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14394_ _14394_/A vssd1 vssd1 vccd1 vccd1 _18476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16133_ _16133_/A vssd1 vssd1 vccd1 vccd1 _19044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13345_ _18641_/Q _13345_/B vssd1 vssd1 vccd1 vccd1 _13345_/X sky130_fd_sc_hd__or2_1
X_10557_ _10557_/A vssd1 vssd1 vccd1 vccd1 _11247_/A sky130_fd_sc_hd__inv_2
XFILLER_155_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09196__A _10622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16064_ _16774_/A vssd1 vssd1 vccd1 vccd1 _16064_/X sky130_fd_sc_hd__clkbuf_1
X_13276_ _13015_/A _13130_/X _12749_/A _18059_/A vssd1 vssd1 vccd1 vccd1 _13276_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10488_ _19254_/Q _19025_/Q _18956_/Q _19350_/Q _10389_/S _09483_/X vssd1 vssd1 vccd1
+ vccd1 _10488_/X sky130_fd_sc_hd__mux4_1
X_15015_ _17751_/A _15015_/B vssd1 vssd1 vccd1 vccd1 _15016_/B sky130_fd_sc_hd__nor2_1
X_12227_ _14568_/A _11966_/B _12173_/Y vssd1 vssd1 vccd1 vccd1 _12227_/X sky130_fd_sc_hd__a21o_1
XFILLER_123_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19823_ _19866_/CLK _19823_/D vssd1 vssd1 vccd1 vccd1 _19823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12158_ _11139_/A _18509_/Q _12328_/A vssd1 vssd1 vccd1 vccd1 _13598_/A sky130_fd_sc_hd__mux2_4
XFILLER_97_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10741__A1 _09629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ _11119_/A _11109_/B vssd1 vssd1 vccd1 vccd1 _11109_/Y sky130_fd_sc_hd__nor2_1
X_19754_ _19755_/CLK _19754_/D vssd1 vssd1 vccd1 vccd1 _19754_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16966_ _16977_/A vssd1 vssd1 vccd1 vccd1 _16975_/S sky130_fd_sc_hd__buf_4
XANTENNA__12350__A _14289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12089_ _12089_/A _12089_/B vssd1 vssd1 vccd1 vccd1 _12096_/B sky130_fd_sc_hd__xor2_4
XFILLER_96_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15680__A1 _15510_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18705_ _19612_/CLK _18705_/D vssd1 vssd1 vccd1 vccd1 _18705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15917_ _15917_/A vssd1 vssd1 vccd1 vccd1 _18960_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14976__S _14997_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19685_ _19689_/CLK _19685_/D vssd1 vssd1 vccd1 vccd1 _19685_/Q sky130_fd_sc_hd__dfxtp_2
X_16897_ _16897_/A vssd1 vssd1 vccd1 vccd1 _19360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17352__S _17352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18636_ _19081_/CLK _18636_/D vssd1 vssd1 vccd1 vccd1 _18636_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15848_ _14918_/X _18930_/Q _15852_/S vssd1 vssd1 vccd1 vccd1 _15849_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18567_ _18567_/CLK _18567_/D vssd1 vssd1 vccd1 vccd1 _18567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15779_ _15779_/A vssd1 vssd1 vccd1 vccd1 _18899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13181__A _18623_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17518_ _19621_/Q _16718_/X _17518_/S vssd1 vssd1 vccd1 vccd1 _17519_/A sky130_fd_sc_hd__mux2_1
X_18498_ _19693_/CLK _18498_/D vssd1 vssd1 vccd1 vccd1 _18498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17449_ _16825_/X _19590_/Q _17457_/S vssd1 vssd1 vccd1 vccd1 _17450_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19119_ _19569_/CLK _19119_/D vssd1 vssd1 vccd1 vccd1 _19119_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_141_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12244__B _12244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17527__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12721__A2 _12742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15671__A1 _15497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09705_ _19429_/Q _19205_/Q _19722_/Q _19173_/Q _09545_/S _10080_/A vssd1 vssd1 vccd1
+ vccd1 _09705_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16667__A _16667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09636_ _10349_/A vssd1 vssd1 vccd1 vccd1 _09636_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_66_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09567_ _19658_/Q _19075_/Q _19112_/Q _18718_/Q _09553_/X _09144_/A vssd1 vssd1 vccd1
+ vccd1 _09568_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10248__B1 _09681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11604__A _13570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09498_ _10650_/S vssd1 vssd1 vccd1 vccd1 _10581_/S sky130_fd_sc_hd__buf_2
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10799__A1 _09409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11996__B1 _17730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17498__A _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10894__S1 _10785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11460_ _11460_/A vssd1 vssd1 vccd1 vccd1 _11460_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10411_ _10412_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _10413_/A sky130_fd_sc_hd__and2_1
XFILLER_99_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11391_ _14801_/A _11391_/B vssd1 vssd1 vccd1 vccd1 _11723_/A sky130_fd_sc_hd__nand2_2
X_13130_ _13130_/A vssd1 vssd1 vccd1 vccd1 _13130_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10342_ _18832_/Q _19386_/Q _19548_/Q _18800_/Q _09734_/A _09610_/A vssd1 vssd1 vccd1
+ vccd1 _10342_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10971__A1 _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13061_ _18330_/Q _13056_/C _13060_/Y vssd1 vssd1 vccd1 vccd1 _18330_/D sky130_fd_sc_hd__o21a_1
XFILLER_3_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10273_ _10266_/X _10268_/X _10270_/X _10272_/X _09248_/A vssd1 vssd1 vccd1 vccd1
+ _10273_/X sky130_fd_sc_hd__a221o_2
XANTENNA__18122__A _19828_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12012_ _11975_/A _14093_/A _11978_/A _11978_/B vssd1 vssd1 vccd1 vccd1 _12013_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input48_A io_ibus_inst[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16820_ _16819_/X _19330_/Q _16823_/S vssd1 vssd1 vccd1 vccd1 _16821_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16751_ _16751_/A vssd1 vssd1 vccd1 vccd1 _19308_/D sky130_fd_sc_hd__clkbuf_1
X_13963_ _13963_/A vssd1 vssd1 vccd1 vccd1 _18431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10487__B1 _10593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15702_ _18865_/Q _15542_/X _15708_/S vssd1 vssd1 vccd1 vccd1 _15703_/A sky130_fd_sc_hd__mux2_1
X_12914_ _18283_/Q vssd1 vssd1 vccd1 vccd1 _12925_/C sky130_fd_sc_hd__clkbuf_1
X_19470_ _19472_/CLK _19470_/D vssd1 vssd1 vccd1 vccd1 _19470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13894_ _13894_/A vssd1 vssd1 vccd1 vccd1 _13931_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16682_ _16682_/A vssd1 vssd1 vccd1 vccd1 _19287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18421_ _18506_/CLK _18421_/D vssd1 vssd1 vccd1 vccd1 _18421_/Q sky130_fd_sc_hd__dfxtp_1
X_12845_ _18263_/Q _12841_/C _12844_/Y vssd1 vssd1 vccd1 vccd1 _18263_/D sky130_fd_sc_hd__o21a_1
X_15633_ _15633_/A vssd1 vssd1 vccd1 vccd1 _18834_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12228__A1 _12493_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11514__A _11514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _18402_/CLK _18352_/D vssd1 vssd1 vccd1 vccd1 _18352_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15564_ _16819_/A vssd1 vssd1 vccd1 vccd1 _15564_/X sky130_fd_sc_hd__clkbuf_2
X_12776_ _19784_/Q _12753_/A _12774_/X _12775_/X vssd1 vssd1 vccd1 vccd1 _12777_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__17167__A1 _13230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11987__A0 _11978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _17303_/A vssd1 vssd1 vccd1 vccd1 _19525_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _18350_/Q _15263_/A vssd1 vssd1 vccd1 vccd1 _11888_/C sky130_fd_sc_hd__and2_1
X_14515_ _18525_/Q _12692_/X _14513_/X _14514_/X vssd1 vssd1 vccd1 vccd1 _18525_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18283_ _19759_/CLK _18283_/D vssd1 vssd1 vccd1 vccd1 _18283_/Q sky130_fd_sc_hd__dfxtp_1
X_15495_ _18786_/Q _15494_/X _15504_/S vssd1 vssd1 vccd1 vccd1 _15496_/A sky130_fd_sc_hd__mux2_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15420__S _15426_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17234_ _17234_/A vssd1 vssd1 vccd1 vccd1 _19496_/D sky130_fd_sc_hd__clkbuf_1
X_11658_ _12152_/B vssd1 vssd1 vccd1 vccd1 _11788_/B sky130_fd_sc_hd__buf_2
X_14446_ _18495_/Q _19733_/Q _14454_/S vssd1 vssd1 vccd1 vccd1 _14447_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11739__A0 _12465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10609_ _10956_/A vssd1 vssd1 vccd1 vccd1 _10830_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17165_ _19476_/Q _17164_/X _17172_/S vssd1 vssd1 vccd1 vccd1 _17166_/A sky130_fd_sc_hd__mux2_1
X_14377_ _14377_/A vssd1 vssd1 vccd1 vccd1 _18470_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10637__S1 _10634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11589_ _11688_/A _11688_/B vssd1 vssd1 vccd1 vccd1 _11618_/A sky130_fd_sc_hd__nand2_2
XFILLER_116_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13328_ _19680_/Q _12668_/X _12768_/X _18404_/Q vssd1 vssd1 vccd1 vccd1 _13329_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_116_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16116_ _16116_/A vssd1 vssd1 vccd1 vccd1 _16129_/S sky130_fd_sc_hd__buf_6
XFILLER_127_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17855__B _19728_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17096_ _17096_/A vssd1 vssd1 vccd1 vccd1 _19448_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13259_ _13217_/X _13248_/Y _13258_/X _13229_/X _18629_/Q vssd1 vssd1 vccd1 vccd1
+ _13259_/X sky130_fd_sc_hd__a32o_4
X_16047_ _16047_/A vssd1 vssd1 vccd1 vccd1 _19017_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16251__S _16257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19806_ _19806_/CLK _19806_/D vssd1 vssd1 vccd1 vccd1 _19806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17998_ _18033_/A _17998_/B _18000_/B vssd1 vssd1 vccd1 vccd1 _19784_/D sky130_fd_sc_hd__nor3_1
XFILLER_38_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19737_ _19738_/CLK _19737_/D vssd1 vssd1 vccd1 vccd1 _19737_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__11408__B _12537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16949_ _16784_/X _19383_/Q _16953_/S vssd1 vssd1 vccd1 vccd1 _16950_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19668_ _19786_/CLK _19668_/D vssd1 vssd1 vccd1 vccd1 _19668_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_65_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10573__S0 _10466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09421_ _09421_/A _09421_/B vssd1 vssd1 vccd1 vccd1 _09421_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18619_ _18623_/CLK _18619_/D vssd1 vssd1 vccd1 vccd1 _18619_/Q sky130_fd_sc_hd__dfxtp_2
X_19599_ _19599_/CLK _19599_/D vssd1 vssd1 vccd1 vccd1 _19599_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11424__A _11821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17810__S _17816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09352_ _09352_/A vssd1 vssd1 vccd1 vccd1 _09353_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_21_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09283_ _09283_/A vssd1 vssd1 vccd1 vccd1 _09284_/A sky130_fd_sc_hd__buf_2
XANTENNA__16426__S _16428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10876__S1 _10616_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18207__A _18207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13195__A2 _13123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10402__A0 _18831_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17765__B _18488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13086__A _18626_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17781__A _17781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10800__S1 _10772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10960_ _10960_/A vssd1 vssd1 vccd1 vccd1 _10960_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10564__S0 _10466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09619_ _10175_/A _09619_/B vssd1 vssd1 vccd1 vccd1 _09619_/Y sky130_fd_sc_hd__nor2_1
X_10891_ _10844_/A _10890_/X _10793_/A vssd1 vssd1 vccd1 vccd1 _10891_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12630_ _18254_/Q _12582_/X _12528_/X _19843_/Q _12629_/X vssd1 vssd1 vccd1 vccd1
+ _12630_/X sky130_fd_sc_hd__a221o_1
XFILLER_34_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12561_ _12810_/A vssd1 vssd1 vccd1 vccd1 _13042_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__16336__S _16340_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10867__S1 _10365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14300_ _14300_/A _14300_/B vssd1 vssd1 vccd1 vccd1 _14300_/Y sky130_fd_sc_hd__nor2_1
X_11512_ _11512_/A _11520_/D vssd1 vssd1 vccd1 vccd1 _11628_/C sky130_fd_sc_hd__or2_2
X_15280_ _15337_/S vssd1 vssd1 vccd1 vccd1 _15289_/S sky130_fd_sc_hd__buf_2
X_12492_ _12492_/A vssd1 vssd1 vccd1 vccd1 _12492_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14231_ _13823_/A _14038_/Y _14230_/X _14115_/X vssd1 vssd1 vccd1 vccd1 _14231_/X
+ sky130_fd_sc_hd__a211o_1
X_11443_ _11432_/X _12688_/C _11822_/B _11723_/B _11442_/Y vssd1 vssd1 vccd1 vccd1
+ _11443_/X sky130_fd_sc_hd__o2111a_1
XFILLER_138_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16860__A _16917_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11197__B2 _11196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14162_ _14162_/A vssd1 vssd1 vccd1 vccd1 _18442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11374_ _11374_/A _11375_/A _11519_/B vssd1 vssd1 vccd1 vccd1 _13583_/A sky130_fd_sc_hd__or3_1
XFILLER_153_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13113_ _17149_/B _13109_/X _13063_/X vssd1 vssd1 vccd1 vccd1 _13113_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_153_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10325_ _10325_/A _10325_/B vssd1 vssd1 vccd1 vccd1 _10325_/Y sky130_fd_sc_hd__nor2_1
X_18970_ _19331_/CLK _18970_/D vssd1 vssd1 vccd1 vccd1 _18970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14093_ _14093_/A _14089_/B vssd1 vssd1 vccd1 vccd1 _14093_/X sky130_fd_sc_hd__or2b_1
XANTENNA__12146__A0 _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17921_ _19817_/Q _19819_/Q _19818_/Q _18089_/A vssd1 vssd1 vccd1 vccd1 _18097_/A
+ sky130_fd_sc_hd__and4_1
X_13044_ _13045_/B _13045_/C _18326_/Q vssd1 vssd1 vccd1 vccd1 _13046_/B sky130_fd_sc_hd__a21oi_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09474__A _10764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10256_ _18602_/Q _19291_/Q _10256_/S vssd1 vssd1 vccd1 vccd1 _10256_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17852_ _17852_/A vssd1 vssd1 vccd1 vccd1 _19726_/D sky130_fd_sc_hd__clkbuf_1
X_10187_ _09867_/A _10184_/Y _10186_/Y _11180_/A vssd1 vssd1 vccd1 vccd1 _10187_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16803_ _16803_/A vssd1 vssd1 vccd1 vccd1 _16803_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13646__A0 _13667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17783_ _17783_/A _17783_/B vssd1 vssd1 vccd1 vccd1 _17840_/A sky130_fd_sc_hd__nand2_8
X_14995_ _16718_/A vssd1 vssd1 vccd1 vccd1 _16822_/A sky130_fd_sc_hd__buf_2
X_19522_ _19818_/CLK _19522_/D vssd1 vssd1 vccd1 vccd1 _19522_/Q sky130_fd_sc_hd__dfxtp_1
X_16734_ _16734_/A vssd1 vssd1 vccd1 vccd1 _16734_/X sky130_fd_sc_hd__clkbuf_2
X_13946_ _13946_/A vssd1 vssd1 vccd1 vccd1 _13946_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19453_ _19714_/CLK _19453_/D vssd1 vssd1 vccd1 vccd1 _19453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16665_ _19282_/Q _16664_/X _16671_/S vssd1 vssd1 vccd1 vccd1 _16666_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13877_ _13742_/X _13746_/X _13877_/S vssd1 vssd1 vccd1 vccd1 _13877_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18404_ _19689_/CLK _18404_/D vssd1 vssd1 vccd1 vccd1 _18404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15616_ _15662_/S vssd1 vssd1 vccd1 vccd1 _15625_/S sky130_fd_sc_hd__buf_2
X_12828_ _12830_/B _12830_/C _12827_/Y vssd1 vssd1 vccd1 vccd1 _18258_/D sky130_fd_sc_hd__o21a_1
X_19384_ _19709_/CLK _19384_/D vssd1 vssd1 vccd1 vccd1 _19384_/Q sky130_fd_sc_hd__dfxtp_1
X_16596_ _16596_/A vssd1 vssd1 vccd1 vccd1 _19253_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10307__S0 _09701_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18335_ _19082_/CLK _18335_/D vssd1 vssd1 vccd1 vccd1 _18335_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15547_ _15547_/A vssd1 vssd1 vccd1 vccd1 _18802_/D sky130_fd_sc_hd__clkbuf_1
X_12759_ _18301_/Q _12758_/X _16211_/B vssd1 vssd1 vccd1 vccd1 _12759_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14555__A _14555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16246__S _16246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15150__S _15153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18266_ _19779_/CLK _18266_/D vssd1 vssd1 vccd1 vccd1 _18266_/Q sky130_fd_sc_hd__dfxtp_1
X_15478_ _15478_/A vssd1 vssd1 vccd1 vccd1 _18780_/D sky130_fd_sc_hd__clkbuf_1
X_17217_ _17217_/A vssd1 vssd1 vccd1 vccd1 _19491_/D sky130_fd_sc_hd__clkbuf_1
X_14429_ _18489_/Q _18521_/Q _15087_/S vssd1 vssd1 vccd1 vccd1 _14430_/A sky130_fd_sc_hd__mux2_1
X_18197_ _18197_/A _18200_/B vssd1 vssd1 vccd1 vccd1 _18197_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_14_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17148_ _17148_/A vssd1 vssd1 vccd1 vccd1 _19471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10935__A1 _10772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15386__A _15397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09970_ _18839_/Q _19393_/Q _19555_/Q _18807_/Q _09803_/A _09881_/A vssd1 vssd1 vccd1
+ vccd1 _09970_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17079_ _17079_/A vssd1 vssd1 vccd1 vccd1 _19440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09384__A _10068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17805__S _17805_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10794__S0 _10934_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13637__A0 _11843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15325__S _15333_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09404_ _09404_/A vssd1 vssd1 vccd1 vccd1 _09940_/A sky130_fd_sc_hd__buf_4
XANTENNA__17540__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09335_ _18977_/Q vssd1 vssd1 vccd1 vccd1 _09336_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10849__S1 _10634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09559__A _10417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ _18530_/Q vssd1 vssd1 vccd1 vccd1 _16212_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_180_clock clkbuf_opt_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19540_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__17776__A _17776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09197_ _11102_/A vssd1 vssd1 vccd1 vccd1 _11097_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16680__A _16680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14117__A1 _12013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10932__S _10932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10110_ _10167_/A _10110_/B vssd1 vssd1 vccd1 vccd1 _10110_/X sky130_fd_sc_hd__or2_1
XANTENNA__14668__A2 _12660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12679__A1 _19662_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11090_ _09695_/A _11087_/X _11089_/X vssd1 vssd1 vccd1 vccd1 _11090_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17067__A0 _16743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10041_ _19522_/Q _19136_/Q _19586_/Q _18742_/Q _09952_/S _10029_/X vssd1 vssd1 vccd1
+ vccd1 _10042_/B sky130_fd_sc_hd__mux4_1
XFILLER_76_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13800_ _14089_/A _13800_/B vssd1 vssd1 vccd1 vccd1 _13800_/X sky130_fd_sc_hd__or2_1
XFILLER_21_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13544__A _13563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17016__A _17062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11992_ _18362_/Q vssd1 vssd1 vccd1 vccd1 _13265_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14780_ input29/X _14703_/A _14779_/X _14732_/X vssd1 vssd1 vccd1 vccd1 _16661_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_63_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10943_ _10950_/A _10938_/X _10942_/X _10728_/X vssd1 vssd1 vccd1 vccd1 _10944_/C
+ sky130_fd_sc_hd__o211a_1
X_13731_ _13783_/B _13590_/X _13728_/X _13730_/X vssd1 vssd1 vccd1 vccd1 _13731_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10311__C1 _09247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_133_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19079_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16450_ _16450_/A vssd1 vssd1 vccd1 vccd1 _19186_/D sky130_fd_sc_hd__clkbuf_1
X_13662_ _12355_/A _13936_/B _13668_/S vssd1 vssd1 vccd1 vccd1 _13662_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10874_ _19506_/Q _19120_/Q _19570_/Q _18726_/Q _10614_/X _10616_/X vssd1 vssd1 vccd1
+ vccd1 _10875_/B sky130_fd_sc_hd__mux4_1
XFILLER_32_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _15401_/A vssd1 vssd1 vccd1 vccd1 _18747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12613_ _18253_/Q _12604_/X _12528_/A _19842_/Q _12612_/X vssd1 vssd1 vccd1 vccd1
+ _12613_/X sky130_fd_sc_hd__a221o_2
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16381_ _16381_/A vssd1 vssd1 vccd1 vccd1 _19156_/D sky130_fd_sc_hd__clkbuf_1
X_13593_ _13737_/A vssd1 vssd1 vccd1 vccd1 _13594_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18120_ _18120_/A _18120_/B _18120_/C vssd1 vssd1 vccd1 vccd1 _19827_/D sky130_fd_sc_hd__nor3_1
X_12544_ _12585_/A vssd1 vssd1 vccd1 vccd1 _13156_/A sky130_fd_sc_hd__buf_2
X_15332_ _15332_/A vssd1 vssd1 vccd1 vccd1 _18717_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_148_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19436_/CLK sky130_fd_sc_hd__clkbuf_16
X_18051_ _19803_/Q _18051_/B _18051_/C vssd1 vssd1 vccd1 vccd1 _18053_/B sky130_fd_sc_hd__and3_1
X_15263_ _15263_/A _15263_/B vssd1 vssd1 vccd1 vccd1 _15263_/X sky130_fd_sc_hd__or2_1
X_12475_ _12475_/A vssd1 vssd1 vccd1 vccd1 _12475_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_126_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17002_ _17002_/A vssd1 vssd1 vccd1 vccd1 _19406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11426_ _12532_/A _12567_/A vssd1 vssd1 vccd1 vccd1 _15241_/A sky130_fd_sc_hd__or2_1
X_14214_ _14216_/A _14216_/B vssd1 vssd1 vccd1 vccd1 _14215_/B sky130_fd_sc_hd__nor2_1
X_15194_ _16696_/A vssd1 vssd1 vccd1 vccd1 _15194_/X sky130_fd_sc_hd__buf_2
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_188_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14145_ _14314_/A _14145_/B vssd1 vssd1 vccd1 vccd1 _14145_/Y sky130_fd_sc_hd__nor2_1
X_11357_ _11375_/A _11640_/A vssd1 vssd1 vccd1 vccd1 _11357_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12119__A0 _14163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10308_ _18832_/Q _19386_/Q _19548_/Q _18800_/Q _09700_/A _10306_/A vssd1 vssd1 vccd1
+ vccd1 _10309_/B sky130_fd_sc_hd__mux4_1
XFILLER_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14076_ _14250_/A _14074_/B _14040_/X _14075_/X vssd1 vssd1 vccd1 vccd1 _14076_/X
+ sky130_fd_sc_hd__o211a_1
X_18953_ _19659_/CLK _18953_/D vssd1 vssd1 vccd1 vccd1 _18953_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output79_A _12066_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11017__S1 _09480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11288_ _11207_/A _11219_/X _11278_/Y _11287_/X vssd1 vssd1 vccd1 vccd1 _11288_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_112_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17904_ _12315_/A _11997_/X _12318_/Y _12321_/X _12802_/X vssd1 vssd1 vccd1 vccd1
+ _19753_/D sky130_fd_sc_hd__a221oi_1
X_13027_ _13035_/D vssd1 vssd1 vccd1 vccd1 _13033_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_140_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10239_ _10239_/A vssd1 vssd1 vccd1 vccd1 _10239_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18884_ _19631_/CLK _18884_/D vssd1 vssd1 vccd1 vccd1 _18884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15608__A1 _15510_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10776__S0 _10724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17835_ _17835_/A vssd1 vssd1 vccd1 vccd1 _19718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17766_ _17765_/A _17765_/C _18488_/Q vssd1 vssd1 vccd1 vccd1 _17766_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_35_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14978_ _17737_/A _14978_/B vssd1 vssd1 vccd1 vccd1 _14980_/B sky130_fd_sc_hd__nor2_1
XFILLER_19_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19505_ _19700_/CLK _19505_/D vssd1 vssd1 vccd1 vccd1 _19505_/Q sky130_fd_sc_hd__dfxtp_1
X_16717_ _16717_/A vssd1 vssd1 vccd1 vccd1 _19298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13929_ _13927_/X _13924_/Y _13928_/X _13795_/A vssd1 vssd1 vccd1 vccd1 _13930_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_62_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17697_ _17701_/A _17701_/C vssd1 vssd1 vccd1 vccd1 _17697_/Y sky130_fd_sc_hd__xnor2_1
X_19436_ _19436_/CLK _19436_/D vssd1 vssd1 vccd1 vccd1 _19436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16648_ _16648_/A vssd1 vssd1 vccd1 vccd1 _16648_/X sky130_fd_sc_hd__buf_2
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19367_ _19625_/CLK _19367_/D vssd1 vssd1 vccd1 vccd1 _19367_/Q sky130_fd_sc_hd__dfxtp_1
X_16579_ _19245_/Q vssd1 vssd1 vccd1 vccd1 _16580_/A sky130_fd_sc_hd__clkbuf_1
X_09120_ _18556_/Q vssd1 vssd1 vccd1 vccd1 _14511_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18318_ _18330_/CLK _18318_/D vssd1 vssd1 vccd1 vccd1 _18318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09379__A _10395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19298_ _19620_/CLK _19298_/D vssd1 vssd1 vccd1 vccd1 _19298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10700__S0 _10886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18249_ _18249_/A _18249_/B _18249_/C vssd1 vssd1 vccd1 vccd1 _19871_/D sky130_fd_sc_hd__nor3_1
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09953_ _09810_/A _09952_/X _10044_/A vssd1 vssd1 vccd1 vccd1 _09953_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_131_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09884_ _09320_/X _09871_/Y _09876_/X _09878_/Y _09883_/Y vssd1 vssd1 vccd1 vccd1
+ _09884_/X sky130_fd_sc_hd__o32a_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_11_0_clock clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_11_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19557_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13389__A2 _13387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_65_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19866_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09318_ _09318_/A vssd1 vssd1 vccd1 vccd1 _09319_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10590_ _19510_/Q _19124_/Q _19574_/Q _18730_/Q _10511_/S _09515_/A vssd1 vssd1 vccd1
+ vccd1 _10591_/B sky130_fd_sc_hd__mux4_1
XFILLER_139_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10072__A1 _09927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14338__A1 _12450_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09249_ _09249_/A vssd1 vssd1 vccd1 vccd1 _09249_/X sky130_fd_sc_hd__buf_4
XANTENNA__10072__B2 _18446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12260_ _09951_/A _12444_/S _12259_/X vssd1 vssd1 vccd1 vccd1 _12286_/A sky130_fd_sc_hd__o21ai_4
XFILLER_154_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11211_ _11475_/A vssd1 vssd1 vccd1 vccd1 _11551_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13539__A _13542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ _12191_/A vssd1 vssd1 vccd1 vccd1 _13529_/B sky130_fd_sc_hd__buf_2
XFILLER_108_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09860__S1 _09841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11142_ _11142_/A vssd1 vssd1 vccd1 vccd1 _11142_/Y sky130_fd_sc_hd__inv_2
Xoutput76 _11978_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[12] sky130_fd_sc_hd__buf_2
XFILLER_89_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput87 _12244_/B vssd1 vssd1 vccd1 vccd1 io_dbus_addr[22] sky130_fd_sc_hd__buf_2
X_15950_ _15076_/X _18976_/Q _15950_/S vssd1 vssd1 vccd1 vccd1 _15951_/A sky130_fd_sc_hd__mux2_1
X_11073_ _10979_/X _11071_/X _11258_/A vssd1 vssd1 vccd1 vccd1 _11073_/X sky130_fd_sc_hd__a21o_1
Xoutput98 _11704_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[3] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10024_ _19618_/Q _19456_/Q _18902_/Q _18672_/Q _10076_/S _09984_/A vssd1 vssd1 vccd1
+ vccd1 _10025_/B sky130_fd_sc_hd__mux4_1
XANTENNA_input30_A io_dbus_rdata[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14901_ _14960_/A vssd1 vssd1 vccd1 vccd1 _14901_/X sky130_fd_sc_hd__buf_2
X_15881_ _15937_/A vssd1 vssd1 vccd1 vccd1 _15950_/S sky130_fd_sc_hd__buf_8
XANTENNA__11875__A2 _11843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17620_ _17620_/A vssd1 vssd1 vccd1 vccd1 _19662_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14832_ _16673_/A vssd1 vssd1 vccd1 vccd1 _16777_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_18_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19595_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17551_ _19635_/Q _16765_/A _17557_/S vssd1 vssd1 vccd1 vccd1 _17552_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14763_ _14763_/A vssd1 vssd1 vccd1 vccd1 _18590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11975_ _11975_/A _12011_/A vssd1 vssd1 vccd1 vccd1 _11978_/A sky130_fd_sc_hd__xor2_4
XANTENNA__17212__A0 _18447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16502_ _16502_/A vssd1 vssd1 vccd1 vccd1 _19210_/D sky130_fd_sc_hd__clkbuf_1
X_13714_ _13796_/A vssd1 vssd1 vccd1 vccd1 _13714_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10926_ _18819_/Q _19373_/Q _19535_/Q _18787_/Q _10668_/A _10906_/A vssd1 vssd1 vccd1
+ vccd1 _10926_/X sky130_fd_sc_hd__mux4_1
X_17482_ _17482_/A vssd1 vssd1 vccd1 vccd1 _19604_/D sky130_fd_sc_hd__clkbuf_1
X_14694_ _14694_/A _14694_/B vssd1 vssd1 vccd1 vccd1 _14695_/A sky130_fd_sc_hd__and2_1
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19221_ _19543_/CLK _19221_/D vssd1 vssd1 vccd1 vccd1 _19221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16433_ _16501_/S vssd1 vssd1 vccd1 vccd1 _16442_/S sky130_fd_sc_hd__buf_2
X_13645_ _13642_/X _13996_/B _13741_/S vssd1 vssd1 vccd1 vccd1 _13811_/A sky130_fd_sc_hd__mux2_1
X_10857_ _10857_/A _10857_/B vssd1 vssd1 vccd1 vccd1 _10857_/X sky130_fd_sc_hd__or2_2
XFILLER_60_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19152_ _19703_/CLK _19152_/D vssd1 vssd1 vccd1 vccd1 _19152_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09199__A _09640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16364_ _16364_/A vssd1 vssd1 vccd1 vccd1 _19148_/D sky130_fd_sc_hd__clkbuf_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13576_ _13657_/S vssd1 vssd1 vccd1 vccd1 _13668_/S sky130_fd_sc_hd__buf_2
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _18590_/Q _19279_/Q _10788_/S vssd1 vssd1 vccd1 vccd1 _10788_/X sky130_fd_sc_hd__mux2_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18103_ _18102_/B _18102_/C _19821_/Q vssd1 vssd1 vccd1 vccd1 _18104_/C sky130_fd_sc_hd__a21oi_1
XFILLER_173_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15315_ _15315_/A vssd1 vssd1 vccd1 vccd1 _18709_/D sky130_fd_sc_hd__clkbuf_1
X_12527_ _12583_/A vssd1 vssd1 vccd1 vccd1 _12528_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19083_ _19632_/CLK _19083_/D vssd1 vssd1 vccd1 vccd1 _19083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16295_ _16295_/A vssd1 vssd1 vccd1 vccd1 _19118_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18034_ _18034_/A vssd1 vssd1 vccd1 vccd1 _18199_/A sky130_fd_sc_hd__clkbuf_4
X_15246_ _18683_/Q _11820_/B _15260_/S vssd1 vssd1 vccd1 vccd1 _15247_/A sky130_fd_sc_hd__mux2_1
X_12458_ _12458_/A _12466_/B vssd1 vssd1 vccd1 vccd1 _12459_/A sky130_fd_sc_hd__and2_2
XFILLER_172_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11409_ _18545_/Q vssd1 vssd1 vccd1 vccd1 _12533_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_141_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12389_ _12385_/X _12388_/Y _12389_/S vssd1 vssd1 vccd1 vccd1 _12389_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15177_ _15177_/A vssd1 vssd1 vccd1 vccd1 _18662_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09851__S1 _09841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14128_ _14142_/A _14128_/B vssd1 vssd1 vccd1 vccd1 _14128_/X sky130_fd_sc_hd__or2_1
XFILLER_141_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17355__S _17363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13304__A2 _13123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15664__A _16744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18936_ _19395_/CLK _18936_/D vssd1 vssd1 vccd1 vccd1 _18936_/Q sky130_fd_sc_hd__dfxtp_1
X_14059_ _14059_/A _14059_/B vssd1 vssd1 vccd1 vccd1 _14059_/X sky130_fd_sc_hd__or2_1
XFILLER_97_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10749__S0 _10669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18867_ _19397_/CLK _18867_/D vssd1 vssd1 vccd1 vccd1 _18867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17818_ _17840_/A vssd1 vssd1 vccd1 vccd1 _17827_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_95_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18798_ _19640_/CLK _18798_/D vssd1 vssd1 vccd1 vccd1 _18798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17749_ _19685_/Q _17748_/X _17772_/S vssd1 vssd1 vccd1 vccd1 _17750_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11141__B_N _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15603__S _15603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10921__S0 _10919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19419_ _19613_/CLK _19419_/D vssd1 vssd1 vccd1 vccd1 _19419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09103_ _18567_/Q vssd1 vssd1 vccd1 vccd1 _11325_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_109_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16434__S _16442_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12263__A _13615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10790__A_N _10887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19691__D _19691_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17265__S _17269_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09936_ _09936_/A vssd1 vssd1 vccd1 vccd1 _09936_/X sky130_fd_sc_hd__clkbuf_4
X_09867_ _09867_/A vssd1 vssd1 vccd1 vccd1 _10029_/A sky130_fd_sc_hd__buf_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09798_ _09992_/A _09798_/B vssd1 vssd1 vccd1 vccd1 _09798_/X sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_136_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _18352_/Q _11719_/B _11726_/B _11759_/X vssd1 vssd1 vccd1 vccd1 _11768_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _10711_/A _18856_/Q vssd1 vssd1 vccd1 vccd1 _10711_/Y sky130_fd_sc_hd__nor2_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15756__A0 _14808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11691_ _13523_/B _14557_/A _15095_/B vssd1 vssd1 vccd1 vccd1 _11692_/C sky130_fd_sc_hd__mux2_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13430_ _12734_/A _18381_/Q _15242_/B _12640_/A vssd1 vssd1 vccd1 vccd1 _13430_/X
+ sky130_fd_sc_hd__a31o_1
X_10642_ _10638_/A _10641_/X _09409_/A vssd1 vssd1 vccd1 vccd1 _10642_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13361_ _13055_/A _12663_/X _12518_/A _18094_/A _13360_/X vssd1 vssd1 vccd1 vccd1
+ _13361_/X sky130_fd_sc_hd__a221o_1
XFILLER_139_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15749__A _15806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10573_ _19606_/Q _19444_/Q _18890_/Q _18660_/Q _10466_/S _10559_/A vssd1 vssd1 vccd1
+ vccd1 _10574_/B sky130_fd_sc_hd__mux4_1
XFILLER_158_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15100_ _18626_/Q _13566_/X _15097_/X _10691_/X vssd1 vssd1 vccd1 vccd1 _18626_/D
+ sky130_fd_sc_hd__a22o_1
X_12312_ _12371_/A _12290_/B _12285_/A vssd1 vssd1 vccd1 vccd1 _12313_/B sky130_fd_sc_hd__a21oi_2
X_13292_ _19806_/Q _12749_/X _13291_/X vssd1 vssd1 vccd1 vccd1 _14873_/D sky130_fd_sc_hd__a21o_1
X_16080_ _16790_/A vssd1 vssd1 vccd1 vccd1 _16080_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12243_ _19750_/Q vssd1 vssd1 vccd1 vccd1 _12246_/A sky130_fd_sc_hd__clkbuf_4
X_15031_ _14999_/X _15025_/X _15028_/X _15030_/X vssd1 vssd1 vccd1 vccd1 _16728_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_142_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12174_ _12489_/C _12226_/A _12172_/Y _12173_/Y vssd1 vssd1 vccd1 vccd1 _14203_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17681__A0 _19673_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ _10442_/A _11124_/X _09681_/X vssd1 vssd1 vccd1 vccd1 _11125_/Y sky130_fd_sc_hd__o21ai_1
X_19770_ _19859_/CLK _19770_/D vssd1 vssd1 vccd1 vccd1 _19770_/Q sky130_fd_sc_hd__dfxtp_1
X_16982_ _16832_/X _19398_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16983_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18721_ _19630_/CLK _18721_/D vssd1 vssd1 vccd1 vccd1 _18721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09482__A _09482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15933_ _14986_/X _18968_/Q _15935_/S vssd1 vssd1 vccd1 vccd1 _15934_/A sky130_fd_sc_hd__mux2_1
X_11056_ _11056_/A _11056_/B vssd1 vssd1 vccd1 vccd1 _11056_/X sky130_fd_sc_hd__or2_1
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10505__C1 _09392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09910__A1 _09217_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10007_ _10007_/A vssd1 vssd1 vccd1 vccd1 _10007_/X sky130_fd_sc_hd__clkbuf_2
X_18652_ _19699_/CLK _18652_/D vssd1 vssd1 vccd1 vccd1 _18652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11517__A _14584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15864_ _15864_/A vssd1 vssd1 vccd1 vccd1 _18937_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14247__A0 _18449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17603_ _19659_/Q _16841_/A _17605_/S vssd1 vssd1 vccd1 vccd1 _17604_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14798__A1 _13228_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14815_ _14815_/A vssd1 vssd1 vccd1 vccd1 _14829_/B sky130_fd_sc_hd__clkbuf_2
X_18583_ _18585_/CLK _18583_/D vssd1 vssd1 vccd1 vccd1 _18583_/Q sky130_fd_sc_hd__dfxtp_1
X_15795_ _15795_/A vssd1 vssd1 vccd1 vccd1 _18906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17534_ _17534_/A vssd1 vssd1 vccd1 vccd1 _19628_/D sky130_fd_sc_hd__clkbuf_1
X_14746_ _15060_/B vssd1 vssd1 vccd1 vccd1 _14981_/S sky130_fd_sc_hd__clkbuf_2
X_11958_ _11956_/X _11957_/Y _12016_/S vssd1 vssd1 vccd1 vccd1 _11958_/X sky130_fd_sc_hd__mux2_1
X_17465_ _17533_/S vssd1 vssd1 vccd1 vccd1 _17474_/S sky130_fd_sc_hd__clkbuf_4
X_10909_ _19691_/Q vssd1 vssd1 vccd1 vccd1 _10909_/X sky130_fd_sc_hd__buf_4
XFILLER_32_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14677_ _14677_/A _14677_/B vssd1 vssd1 vccd1 vccd1 _14678_/A sky130_fd_sc_hd__and2_1
X_11889_ _17221_/A _11962_/D vssd1 vssd1 vccd1 vccd1 _11889_/Y sky130_fd_sc_hd__nor2_1
X_19204_ _19721_/CLK _19204_/D vssd1 vssd1 vccd1 vccd1 _19204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16416_ _19172_/Q _15570_/X _16424_/S vssd1 vssd1 vccd1 vccd1 _16417_/A sky130_fd_sc_hd__mux2_1
X_13628_ _13650_/A vssd1 vssd1 vccd1 vccd1 _13991_/S sky130_fd_sc_hd__clkbuf_2
X_17396_ _16749_/X _19566_/Q _17402_/S vssd1 vssd1 vccd1 vccd1 _17397_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09426__B1 _09425_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12067__B _12067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09977__A1 _10010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19135_ _19716_/CLK _19135_/D vssd1 vssd1 vccd1 vccd1 _19135_/Q sky130_fd_sc_hd__dfxtp_1
X_16347_ _16122_/X _19142_/Q _16351_/S vssd1 vssd1 vccd1 vccd1 _16348_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14970__A1 _13345_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13559_ _09094_/A _13536_/X _13537_/A _18424_/Q vssd1 vssd1 vccd1 vccd1 _13560_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18035__A _18199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19066_ _19810_/CLK _19066_/D vssd1 vssd1 vccd1 vccd1 _19066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16278_ _16278_/A vssd1 vssd1 vccd1 vccd1 _19111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18017_ _19791_/Q _18015_/B _17993_/X vssd1 vssd1 vccd1 vccd1 _18017_/Y sky130_fd_sc_hd__a21oi_1
X_15229_ _16731_/A vssd1 vssd1 vccd1 vccd1 _15229_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09392__A _09392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09721_ _11186_/S vssd1 vssd1 vccd1 vccd1 _09721_/X sky130_fd_sc_hd__buf_4
XFILLER_80_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18919_ _19541_/CLK _18919_/D vssd1 vssd1 vccd1 vccd1 _18919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17424__A0 _16790_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10198__S1 _09978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09652_ _19624_/Q _19462_/Q _18908_/Q _18678_/Q _09700_/A _09636_/X vssd1 vssd1 vccd1
+ vccd1 _09652_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10331__A _10331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14789__A1 _14788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09583_ _09583_/A vssd1 vssd1 vccd1 vccd1 _10328_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14644__A1_N input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15333__S _15333_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11162__A _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__S1 _10368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16164__S _16172_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14961__A1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18152__A1 _19837_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10578__A2 _10568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_62_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17784__A _17840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09815__S1 _09810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09919_ _09919_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _09919_/X sky130_fd_sc_hd__or2_1
XFILLER_101_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12930_ _18287_/Q _18286_/Q _12930_/C _12930_/D vssd1 vssd1 vccd1 vccd1 _12932_/B
+ sky130_fd_sc_hd__and4_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _12991_/A vssd1 vssd1 vccd1 vccd1 _12904_/A sky130_fd_sc_hd__buf_2
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14648__A _14648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _14612_/A _14600_/B vssd1 vssd1 vccd1 vccd1 _18555_/D sky130_fd_sc_hd__nand2_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11812_ _11783_/B _11787_/B _11811_/Y vssd1 vssd1 vccd1 vccd1 _11813_/B sky130_fd_sc_hd__o21a_1
X_15580_ _16835_/A vssd1 vssd1 vccd1 vccd1 _15580_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _11822_/B _15241_/B _12790_/X _12791_/X vssd1 vssd1 vccd1 vccd1 _18205_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _15134_/A vssd1 vssd1 vccd1 vccd1 _16919_/C sky130_fd_sc_hd__clkbuf_4
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11785_/A _11784_/A vssd1 vssd1 vccd1 vccd1 _11745_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10387__S _10387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17250_ _19501_/Q _16639_/X _17258_/S vssd1 vssd1 vccd1 vccd1 _17251_/A sky130_fd_sc_hd__mux2_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _14462_/A vssd1 vssd1 vccd1 vccd1 _18502_/D sky130_fd_sc_hd__clkbuf_1
X_11674_ _18344_/Q _18337_/Q _11673_/Y _18339_/Q _18346_/Q vssd1 vssd1 vccd1 vccd1
+ _11674_/X sky130_fd_sc_hd__a32o_1
XFILLER_30_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16201_ _16122_/X _19073_/Q _16205_/S vssd1 vssd1 vccd1 vccd1 _16202_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13413_ _18379_/Q _13413_/B vssd1 vssd1 vccd1 vccd1 _13413_/X sky130_fd_sc_hd__or2_1
X_17181_ _18438_/Q _12727_/X _17184_/S vssd1 vssd1 vccd1 vccd1 _17181_/X sky130_fd_sc_hd__mux2_1
X_10625_ _18825_/Q _19379_/Q _19541_/Q _18793_/Q _10353_/A _10548_/X vssd1 vssd1 vccd1
+ vccd1 _10625_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14393_ _17701_/B _18508_/Q _14395_/S vssd1 vssd1 vccd1 vccd1 _14394_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10113__S1 _10103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09477__A _09522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16132_ _16131_/X _19044_/Q _16135_/S vssd1 vssd1 vccd1 vccd1 _16133_/A sky130_fd_sc_hd__mux2_1
X_13344_ _19491_/Q _13203_/X _13338_/X _13339_/X _13343_/X vssd1 vssd1 vccd1 vccd1
+ _13345_/B sky130_fd_sc_hd__a2111o_2
X_10556_ _11081_/A _10556_/B vssd1 vssd1 vccd1 vccd1 _10557_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12615__B _12615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16063_ _16063_/A vssd1 vssd1 vccd1 vccd1 _19022_/D sky130_fd_sc_hd__clkbuf_1
X_13275_ _19805_/Q vssd1 vssd1 vccd1 vccd1 _18059_/A sky130_fd_sc_hd__clkbuf_2
X_10487_ _09501_/A _10486_/X _10593_/A vssd1 vssd1 vccd1 vccd1 _10487_/X sky130_fd_sc_hd__a21o_1
XFILLER_136_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15014_ _18484_/Q _15015_/B vssd1 vssd1 vccd1 vccd1 _15037_/C sky130_fd_sc_hd__and2_1
XFILLER_142_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12226_ _12226_/A vssd1 vssd1 vccd1 vccd1 _12345_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_170_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15418__S _15426_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19822_ _19822_/CLK _19822_/D vssd1 vssd1 vccd1 vccd1 _19822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12157_ _14192_/A _12157_/B vssd1 vssd1 vccd1 vccd1 _12160_/A sky130_fd_sc_hd__xnor2_1
XFILLER_68_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11108_ _18766_/Q _18995_/Q _18926_/Q _19224_/Q _10279_/S _10390_/A vssd1 vssd1 vccd1
+ vccd1 _11109_/B sky130_fd_sc_hd__mux4_1
X_19753_ _19753_/CLK _19753_/D vssd1 vssd1 vccd1 vccd1 _19753_/Q sky130_fd_sc_hd__dfxtp_4
X_16965_ _16965_/A vssd1 vssd1 vccd1 vccd1 _19390_/D sky130_fd_sc_hd__clkbuf_1
X_12088_ _12040_/A _12040_/B _12066_/A _12087_/X vssd1 vssd1 vccd1 vccd1 _12089_/B
+ sky130_fd_sc_hd__a31o_2
X_11039_ _10973_/A _11038_/X _09208_/A vssd1 vssd1 vccd1 vccd1 _11039_/Y sky130_fd_sc_hd__o21ai_1
X_18704_ _19714_/CLK _18704_/D vssd1 vssd1 vccd1 vccd1 _18704_/Q sky130_fd_sc_hd__dfxtp_1
X_15916_ _14889_/X _18960_/Q _15924_/S vssd1 vssd1 vccd1 vccd1 _15917_/A sky130_fd_sc_hd__mux2_1
X_19684_ _19686_/CLK _19684_/D vssd1 vssd1 vccd1 vccd1 _19684_/Q sky130_fd_sc_hd__dfxtp_2
X_16896_ _19360_/Q _16709_/X _16902_/S vssd1 vssd1 vccd1 vccd1 _16897_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09940__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18635_ _19081_/CLK _18635_/D vssd1 vssd1 vccd1 vccd1 _18635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15847_ _15847_/A vssd1 vssd1 vccd1 vccd1 _18929_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16249__S _16257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15153__S _15153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18566_ _18567_/CLK _18566_/D vssd1 vssd1 vccd1 vccd1 _18566_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09647__B1 _09133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15778_ _14929_/X _18899_/Q _15780_/S vssd1 vssd1 vccd1 vccd1 _15779_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17517_ _17517_/A vssd1 vssd1 vccd1 vccd1 _19620_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13181__B _13181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__S0 _09734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14729_ _16749_/A vssd1 vssd1 vccd1 vccd1 _14729_/X sky130_fd_sc_hd__clkbuf_2
X_18497_ _19693_/CLK _18497_/D vssd1 vssd1 vccd1 vccd1 _18497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17448_ _17448_/A vssd1 vssd1 vccd1 vccd1 _17457_/S sky130_fd_sc_hd__buf_4
XFILLER_21_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17379_ _16829_/X _19559_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _17380_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12806__A _12991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10104__S1 _10103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12954__B1 _12948_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19118_ _19632_/CLK _19118_/D vssd1 vssd1 vccd1 vccd1 _19118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17808__S _17816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19049_ _19632_/CLK _19049_/D vssd1 vssd1 vccd1 vccd1 _19049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15120__B2 _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09704_ _09704_/A vssd1 vssd1 vccd1 vccd1 _10080_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13682__A1 _14045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09635_ _09635_/A vssd1 vssd1 vccd1 vccd1 _10349_/A sky130_fd_sc_hd__buf_2
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10996__A _10996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09566_ _10313_/A _09566_/B vssd1 vssd1 vccd1 vccd1 _09566_/X sky130_fd_sc_hd__or2_1
XFILLER_71_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10248__A1 _10395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11604__B _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09497_ _10631_/A vssd1 vssd1 vccd1 vccd1 _10650_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16683__A _16683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18125__A1 _19828_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10410_ _18440_/Q _09308_/A _09429_/A _10409_/X vssd1 vssd1 vccd1 vccd1 _12482_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11390_ _14900_/A _18427_/Q _14900_/B _18426_/Q vssd1 vssd1 vccd1 vccd1 _11391_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_109_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10420__A1 _09642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10341_ _11185_/A _10341_/B vssd1 vssd1 vccd1 vccd1 _10341_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10236__A _10447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13060_ _17948_/A _13067_/C vssd1 vssd1 vccd1 vccd1 _13060_/Y sky130_fd_sc_hd__nor2_1
X_10272_ _09995_/A _10271_/X _09988_/A vssd1 vssd1 vccd1 vccd1 _10272_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17636__A0 _13212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12011_ _12011_/A vssd1 vssd1 vccd1 vccd1 _14093_/A sky130_fd_sc_hd__buf_2
XFILLER_105_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12451__A _19759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17453__S _17457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16750_ _16749_/X _19308_/Q _16759_/S vssd1 vssd1 vccd1 vccd1 _16751_/A sky130_fd_sc_hd__mux2_1
X_13962_ _18431_/Q _13961_/X _14032_/S vssd1 vssd1 vccd1 vccd1 _13963_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09760__A _10075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15701_ _15701_/A vssd1 vssd1 vccd1 vccd1 _18864_/D sky130_fd_sc_hd__clkbuf_1
X_12913_ _18282_/Q _12908_/B _12912_/Y vssd1 vssd1 vccd1 vccd1 _18282_/D sky130_fd_sc_hd__o21a_1
XFILLER_58_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16681_ _19287_/Q _16680_/X _16687_/S vssd1 vssd1 vccd1 vccd1 _16682_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16069__S _16081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13893_ _13893_/A vssd1 vssd1 vccd1 vccd1 _13894_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18420_ _18509_/CLK _18420_/D vssd1 vssd1 vccd1 vccd1 _18420_/Q sky130_fd_sc_hd__dfxtp_1
X_15632_ _18834_/Q _15545_/X _15636_/S vssd1 vssd1 vccd1 vccd1 _15633_/A sky130_fd_sc_hd__mux2_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _12844_/A _12850_/C vssd1 vssd1 vccd1 vccd1 _12844_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _18386_/CLK _18351_/D vssd1 vssd1 vccd1 vccd1 _18351_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09724__S0 _09721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _15563_/A vssd1 vssd1 vccd1 vccd1 _18807_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _18259_/Q _12604_/A _12748_/A _19816_/Q vssd1 vssd1 vccd1 vccd1 _12775_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _19525_/Q _16718_/X _17302_/S vssd1 vssd1 vccd1 vccd1 _17303_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _14514_/A vssd1 vssd1 vccd1 vccd1 _14514_/X sky130_fd_sc_hd__buf_2
XFILLER_30_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ _18298_/CLK _18282_/D vssd1 vssd1 vccd1 vccd1 _18282_/Q sky130_fd_sc_hd__dfxtp_2
X_11726_ _11726_/A _11726_/B vssd1 vssd1 vccd1 vccd1 _11726_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15494_ _16749_/A vssd1 vssd1 vccd1 vccd1 _15494_/X sky130_fd_sc_hd__buf_2
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17233_ _19496_/Q _17232_/X _17239_/S vssd1 vssd1 vccd1 vccd1 _17234_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14445_ _14502_/S vssd1 vssd1 vccd1 vccd1 _14454_/S sky130_fd_sc_hd__clkbuf_2
X_11657_ _11999_/A vssd1 vssd1 vccd1 vccd1 _12152_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_30_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12936__B1 _17895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17164_ _18433_/Q _13088_/A _17167_/S vssd1 vssd1 vccd1 vccd1 _17164_/X sky130_fd_sc_hd__mux2_1
X_10608_ _10923_/A vssd1 vssd1 vccd1 vccd1 _10956_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14376_ _14861_/A _18502_/Q _14381_/S vssd1 vssd1 vccd1 vccd1 _14377_/A sky130_fd_sc_hd__mux2_1
X_11588_ _12458_/A _11831_/A vssd1 vssd1 vccd1 vccd1 _11688_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16115_ _16825_/A vssd1 vssd1 vccd1 vccd1 _16115_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13327_ _19490_/Q _13235_/X _13236_/X _18371_/Q _13326_/X vssd1 vssd1 vccd1 vccd1
+ _13329_/A sky130_fd_sc_hd__a221o_1
XANTENNA__17628__S _17628_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10539_ _10566_/A _10539_/B vssd1 vssd1 vccd1 vccd1 _10539_/X sky130_fd_sc_hd__or2_1
X_17095_ _16787_/X _19448_/Q _17097_/S vssd1 vssd1 vccd1 vccd1 _17096_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09935__A _10132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16046_ _16045_/X _19017_/Q _16049_/S vssd1 vssd1 vccd1 vccd1 _16047_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14153__A2 _14155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13258_ _18629_/Q _14824_/B _14824_/C _14824_/D vssd1 vssd1 vccd1 vccd1 _13258_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12209_ _12209_/A _14216_/B vssd1 vssd1 vccd1 vccd1 _12237_/A sky130_fd_sc_hd__and2_1
XANTENNA__12361__A _12361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13189_ _18272_/Q _13326_/B _13127_/A _18355_/Q vssd1 vssd1 vccd1 vccd1 _13189_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19805_ _19806_/CLK _19805_/D vssd1 vssd1 vccd1 vccd1 _19805_/Q sky130_fd_sc_hd__dfxtp_1
X_17997_ _19784_/Q _19783_/Q _17997_/C vssd1 vssd1 vccd1 vccd1 _18000_/B sky130_fd_sc_hd__and3_1
XANTENNA__14987__S _14997_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13113__B1 _13063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17363__S _17363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16850__A1 _16639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19736_ _19738_/CLK _19736_/D vssd1 vssd1 vccd1 vccd1 _19736_/Q sky130_fd_sc_hd__dfxtp_1
X_16948_ _16948_/A vssd1 vssd1 vccd1 vccd1 _19382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19667_ _19786_/CLK _19667_/D vssd1 vssd1 vccd1 vccd1 _19667_/Q sky130_fd_sc_hd__dfxtp_4
X_16879_ _16879_/A vssd1 vssd1 vccd1 vccd1 _19352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_10_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09420_ _19532_/Q _19146_/Q _19596_/Q _18752_/Q _09369_/S _09370_/A vssd1 vssd1 vccd1
+ vccd1 _09421_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10573__S1 _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18618_ _18618_/CLK input72/X vssd1 vssd1 vccd1 vccd1 _18618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19598_ _19598_/CLK _19598_/D vssd1 vssd1 vccd1 vccd1 _19598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09715__S0 _09545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09351_ _10712_/A vssd1 vssd1 vccd1 vccd1 _09352_/A sky130_fd_sc_hd__buf_4
X_18549_ _19481_/CLK _18549_/D vssd1 vssd1 vccd1 vccd1 _18549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16707__S _16719_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14717__C_N _15134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15169__A1 _15168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09282_ _09282_/A vssd1 vssd1 vccd1 vccd1 _09283_/A sky130_fd_sc_hd__buf_2
XANTENNA__09191__S1 _09149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12324__A1_N _14578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13719__A2 _12510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14916__A1 _14711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17538__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16442__S _16442_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13086__B _13086_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10261__S0 _09793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09618_ _18846_/Q _19400_/Q _19562_/Q _18814_/Q _10131_/S _09610_/X vssd1 vssd1 vccd1
+ vccd1 _09619_/B sky130_fd_sc_hd__mux4_1
X_10890_ _18755_/Q _18984_/Q _18915_/Q _19213_/Q _11050_/S _09512_/A vssd1 vssd1 vccd1
+ vccd1 _10890_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09706__S0 _09692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09549_ _09549_/A vssd1 vssd1 vccd1 vccd1 _10475_/A sky130_fd_sc_hd__buf_2
XFILLER_24_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12560_ input72/X vssd1 vssd1 vccd1 vccd1 _12810_/A sky130_fd_sc_hd__buf_2
XFILLER_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ _11511_/A _11550_/B _11511_/C vssd1 vssd1 vccd1 vccd1 _11520_/D sky130_fd_sc_hd__or3_1
XFILLER_156_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12446__A _14332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12491_ _12495_/A _12495_/B _12491_/C vssd1 vssd1 vccd1 vccd1 _12492_/A sky130_fd_sc_hd__and3_1
XFILLER_138_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14230_ _14037_/X _14036_/X _14229_/Y _13594_/A vssd1 vssd1 vccd1 vccd1 _14230_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11442_ _18416_/Q vssd1 vssd1 vccd1 vccd1 _11442_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10929__C1 _10821_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14161_ _18442_/Q _14160_/X _14209_/S vssd1 vssd1 vccd1 vccd1 _14162_/A sky130_fd_sc_hd__mux2_1
X_11373_ _18584_/Q _11475_/A _11333_/X _11362_/A _11640_/A vssd1 vssd1 vccd1 vccd1
+ _11481_/B sky130_fd_sc_hd__a2111o_1
XFILLER_166_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14661__A _14677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13112_ _13112_/A vssd1 vssd1 vccd1 vccd1 _17149_/B sky130_fd_sc_hd__clkinv_2
XANTENNA_input60_A io_ibus_inst[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10324_ _18768_/Q _18997_/Q _18928_/Q _19226_/Q _09734_/A _09610_/A vssd1 vssd1 vccd1
+ vccd1 _10325_/B sky130_fd_sc_hd__mux4_1
XFILLER_166_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14092_ _14092_/A _14092_/B vssd1 vssd1 vccd1 vccd1 _14092_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13043_ _18085_/A vssd1 vssd1 vccd1 vccd1 _17935_/A sky130_fd_sc_hd__clkbuf_2
X_17920_ _19815_/Q _19814_/Q _19816_/Q _18079_/A vssd1 vssd1 vccd1 vccd1 _18089_/A
+ sky130_fd_sc_hd__and4_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ _10270_/A _10255_/B vssd1 vssd1 vccd1 vccd1 _10255_/X sky130_fd_sc_hd__or2_1
XFILLER_106_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17851_ _15235_/X _19726_/Q _17853_/S vssd1 vssd1 vccd1 vccd1 _17852_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10186_ _10186_/A _10186_/B vssd1 vssd1 vccd1 vccd1 _10186_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16802_ _16802_/A vssd1 vssd1 vccd1 vccd1 _19324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17782_ _17782_/A vssd1 vssd1 vccd1 vccd1 _19695_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13646__A1 _12381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14994_ _14994_/A _14994_/B vssd1 vssd1 vccd1 vccd1 _16718_/A sky130_fd_sc_hd__and2_4
XFILLER_115_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19521_ _19716_/CLK _19521_/D vssd1 vssd1 vccd1 vccd1 _19521_/Q sky130_fd_sc_hd__dfxtp_1
X_16733_ _16733_/A vssd1 vssd1 vccd1 vccd1 _19303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09945__S0 _09809_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13945_ _14278_/A vssd1 vssd1 vccd1 vccd1 _13949_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13724__B _13724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_184_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19452_ _19452_/CLK _19452_/D vssd1 vssd1 vccd1 vccd1 _19452_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11525__A _13578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16664_ _16664_/A vssd1 vssd1 vccd1 vccd1 _16664_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13876_ _13741_/X _13755_/X _13879_/S vssd1 vssd1 vccd1 vccd1 _13876_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18403_ _19788_/CLK _18403_/D vssd1 vssd1 vccd1 vccd1 _18403_/Q sky130_fd_sc_hd__dfxtp_1
X_15615_ _15615_/A vssd1 vssd1 vccd1 vccd1 _18826_/D sky130_fd_sc_hd__clkbuf_1
X_12827_ _12830_/B _12830_/C _12817_/X vssd1 vssd1 vccd1 vccd1 _12827_/Y sky130_fd_sc_hd__a21oi_1
X_19383_ _19609_/CLK _19383_/D vssd1 vssd1 vccd1 vccd1 _19383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16595_ _19253_/Q vssd1 vssd1 vccd1 vccd1 _16596_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__10880__B2 _10879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10307__S1 _10306_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18334_ _19866_/CLK _18334_/D vssd1 vssd1 vccd1 vccd1 _18334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15546_ _18802_/Q _15545_/X _15552_/S vssd1 vssd1 vccd1 vccd1 _15547_/A sky130_fd_sc_hd__mux2_1
X_12758_ _12732_/X _12757_/X _12780_/S vssd1 vssd1 vccd1 vccd1 _12758_/X sky130_fd_sc_hd__mux2_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18265_ _19779_/CLK _18265_/D vssd1 vssd1 vccd1 vccd1 _18265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11709_ _11704_/Y _11707_/X _12389_/S vssd1 vssd1 vccd1 vccd1 _11709_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15477_ _18780_/Q _15226_/X _15481_/S vssd1 vssd1 vccd1 vccd1 _15478_/A sky130_fd_sc_hd__mux2_1
X_12689_ _18341_/Q _12687_/X _16211_/B vssd1 vssd1 vccd1 vccd1 _12689_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17216_ _19491_/Q _17215_/X _17223_/S vssd1 vssd1 vccd1 vccd1 _17217_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14428_ _14428_/A vssd1 vssd1 vccd1 vccd1 _18488_/D sky130_fd_sc_hd__clkbuf_1
X_18196_ _19853_/Q _19852_/Q _18196_/C vssd1 vssd1 vccd1 vccd1 _18200_/B sky130_fd_sc_hd__and3_1
XFILLER_129_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17147_ _19471_/Q _17146_/X _17155_/S vssd1 vssd1 vccd1 vccd1 _17148_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09786__C1 _09854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16262__S _16268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09250__A1 _09217_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14359_ _14786_/A _18496_/Q _14367_/S vssd1 vssd1 vccd1 vccd1 _14360_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17078_ _16761_/X _19440_/Q _17086_/S vssd1 vssd1 vccd1 vccd1 _17079_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10491__S0 _09522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17882__A _17882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16029_ _15066_/X _19012_/Q _16031_/S vssd1 vssd1 vccd1 vccd1 _16030_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11896__A0 _10601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15087__A0 _18621_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17093__S _17097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10794__S1 _10785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13098__C1 _14612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13637__A1 _12307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19719_ _19720_/CLK _19719_/D vssd1 vssd1 vccd1 vccd1 _19719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09710__C1 _09134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17821__S _17827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09403_ _09403_/A vssd1 vssd1 vccd1 vccd1 _09404_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_111_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13650__A _13650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09334_ _09819_/A vssd1 vssd1 vccd1 vccd1 _09421_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10084__C1 _09135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12793__B_N _13532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09265_ _18571_/Q _18531_/Q vssd1 vssd1 vccd1 vccd1 _09265_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_14_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09196_ _10622_/A vssd1 vssd1 vccd1 vccd1 _11102_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12376__B2 _12502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09241__A1 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16172__S _16172_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13097__A _17781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16900__S _16902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12679__A2 _12668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10040_ _09892_/X _10035_/X _10037_/X _10039_/X _09404_/A vssd1 vssd1 vccd1 vccd1
+ _10040_/X sky130_fd_sc_hd__a221o_2
XFILLER_88_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11991_ _11980_/X _11987_/X _11990_/X vssd1 vssd1 vccd1 vccd1 _11991_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13730_ _14102_/A vssd1 vssd1 vccd1 vccd1 _13730_/X sky130_fd_sc_hd__clkbuf_2
X_10942_ _11060_/A _10942_/B vssd1 vssd1 vccd1 vccd1 _10942_/X sky130_fd_sc_hd__or2_1
XFILLER_44_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13661_ _14289_/B _13925_/B _13668_/S vssd1 vssd1 vccd1 vccd1 _13661_/X sky130_fd_sc_hd__mux2_1
X_10873_ _10873_/A _10873_/B vssd1 vssd1 vccd1 vccd1 _10873_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16347__S _16351_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15251__S _17143_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15400_ _18747_/Q _15223_/X _15406_/S vssd1 vssd1 vccd1 vccd1 _15401_/A sky130_fd_sc_hd__mux2_1
X_12612_ _19778_/Q _12611_/X _12628_/A vssd1 vssd1 vccd1 vccd1 _12612_/X sky130_fd_sc_hd__mux2_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16380_ _19156_/Q _15519_/X _16380_/S vssd1 vssd1 vccd1 vccd1 _16381_/A sky130_fd_sc_hd__mux2_1
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _13729_/B _13724_/B vssd1 vssd1 vccd1 vccd1 _13737_/A sky130_fd_sc_hd__nand2_1
XFILLER_169_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15331_ _18717_/Q _15229_/X _15333_/S vssd1 vssd1 vccd1 vccd1 _15332_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12543_ _18347_/Q _12643_/A _12742_/A _18399_/Q _12542_/X vssd1 vssd1 vccd1 vccd1
+ _12543_/X sky130_fd_sc_hd__a221o_1
XFILLER_129_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12176__A _14203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16871__A _16917_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18050_ _18051_/B _18051_/C _18049_/Y vssd1 vssd1 vccd1 vccd1 _19802_/D sky130_fd_sc_hd__o21a_1
X_15262_ _15262_/A _15262_/B vssd1 vssd1 vccd1 vccd1 _15263_/B sky130_fd_sc_hd__nor2_1
XANTENNA__16750__A0 _16749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12474_ _12472_/A _12474_/B vssd1 vssd1 vccd1 vccd1 _12475_/A sky130_fd_sc_hd__and2b_1
XFILLER_138_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17001_ _19406_/Q _16651_/X _17003_/S vssd1 vssd1 vccd1 vccd1 _17002_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14213_ _14212_/A _13623_/Y _13797_/X _14212_/Y vssd1 vssd1 vccd1 vccd1 _14213_/X
+ sky130_fd_sc_hd__o211a_1
X_11425_ _12530_/A _12686_/A _12519_/A vssd1 vssd1 vccd1 vccd1 _12567_/A sky130_fd_sc_hd__nor3_1
XFILLER_137_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10378__A0 _18831_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09232__A1 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15193_ _15193_/A vssd1 vssd1 vccd1 vccd1 _18667_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12904__A _12904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11052__A_N _10713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14144_ _13970_/S _13656_/X _13899_/X vssd1 vssd1 vccd1 vccd1 _14145_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__15305__A1 _15191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11356_ _11356_/A vssd1 vssd1 vccd1 vccd1 _11356_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10307_ _19612_/Q _19450_/Q _18896_/Q _18666_/Q _09701_/S _10306_/X vssd1 vssd1 vccd1
+ vccd1 _10307_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14075_ _14178_/A _14075_/B vssd1 vssd1 vccd1 vccd1 _14075_/X sky130_fd_sc_hd__or2_1
X_18952_ _19506_/CLK _18952_/D vssd1 vssd1 vccd1 vccd1 _18952_/Q sky130_fd_sc_hd__dfxtp_1
X_11287_ _11337_/A _11528_/A _11358_/B _11299_/A vssd1 vssd1 vccd1 vccd1 _11287_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_140_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17903_ _17902_/Y _11997_/X _12296_/Y _12300_/X _12802_/X vssd1 vssd1 vccd1 vccd1
+ _19752_/D sky130_fd_sc_hd__a221oi_1
X_13026_ _18320_/Q _18319_/Q _18321_/Q _13026_/D vssd1 vssd1 vccd1 vccd1 _13035_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__10225__S0 _10224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10238_ _10238_/A vssd1 vssd1 vccd1 vccd1 _10239_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18883_ _19698_/CLK _18883_/D vssd1 vssd1 vccd1 vccd1 _18883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15426__S _15426_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10776__S1 _10713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17834_ _15210_/X _19718_/Q _17838_/S vssd1 vssd1 vccd1 vccd1 _17835_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10169_ _10093_/A _10168_/X _09230_/A vssd1 vssd1 vccd1 vccd1 _10169_/X sky130_fd_sc_hd__o21a_1
XFILLER_120_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09918__S0 _09914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14977_ _14977_/A vssd1 vssd1 vccd1 vccd1 _18608_/D sky130_fd_sc_hd__clkbuf_1
X_17765_ _17765_/A _18488_/Q _17765_/C vssd1 vssd1 vccd1 vccd1 _17770_/B sky130_fd_sc_hd__or3_1
XFILLER_54_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19504_ _19632_/CLK _19504_/D vssd1 vssd1 vccd1 vccd1 _19504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16716_ _19298_/Q _16715_/X _16719_/S vssd1 vssd1 vccd1 vccd1 _16717_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13928_ _11602_/Y _13891_/A _13925_/B _14089_/A _13797_/A vssd1 vssd1 vccd1 vccd1
+ _13928_/X sky130_fd_sc_hd__o221a_1
XFILLER_75_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17696_ _17696_/A vssd1 vssd1 vccd1 vccd1 _19675_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16647_ _16647_/A vssd1 vssd1 vccd1 vccd1 _19276_/D sky130_fd_sc_hd__clkbuf_1
X_19435_ _19436_/CLK _19435_/D vssd1 vssd1 vccd1 vccd1 _19435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13859_ _14320_/A _13665_/X _14092_/A _13858_/Y vssd1 vssd1 vccd1 vccd1 _13862_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16257__S _16257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16578_ _16578_/A vssd1 vssd1 vccd1 vccd1 _19244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19366_ _19723_/CLK _19366_/D vssd1 vssd1 vccd1 vccd1 _19366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14285__B _14289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18317_ _18329_/CLK _18317_/D vssd1 vssd1 vccd1 vccd1 _18317_/Q sky130_fd_sc_hd__dfxtp_1
X_15529_ _16784_/A vssd1 vssd1 vccd1 vccd1 _15529_/X sky130_fd_sc_hd__clkbuf_2
X_19297_ _19587_/CLK _19297_/D vssd1 vssd1 vccd1 vccd1 _19297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09471__B2 _18456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10700__S1 _09352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18248_ _18247_/B _18247_/C _19871_/Q vssd1 vssd1 vccd1 vccd1 _18249_/C sky130_fd_sc_hd__a21oi_1
XFILLER_136_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15397__A _15397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18179_ _19846_/Q _18177_/B _18178_/Y vssd1 vssd1 vccd1 vccd1 _19846_/D sky130_fd_sc_hd__o21a_1
XANTENNA__14505__S _14565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09395__A _09395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11030__A1 _10548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17816__S _17816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09952_ _18608_/Q _19297_/Q _09952_/S vssd1 vssd1 vccd1 vccd1 _09952_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09883_ _09944_/A _09882_/X _09320_/A vssd1 vssd1 vccd1 vccd1 _09883_/Y sky130_fd_sc_hd__o21ai_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10519__S1 _10238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12294__A0 _12290_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11192__S1 _10329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09317_ _09317_/A vssd1 vssd1 vccd1 vccd1 _09318_/A sky130_fd_sc_hd__buf_2
XFILLER_51_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09248_ _09248_/A vssd1 vssd1 vccd1 vccd1 _09249_/A sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_132_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09179_ _09179_/A vssd1 vssd1 vccd1 vccd1 _09451_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11021__A1 _09407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ _11376_/A vssd1 vssd1 vccd1 vccd1 _11475_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12190_ _12185_/X _12188_/Y _12452_/S vssd1 vssd1 vccd1 vccd1 _12190_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11141_ _12491_/C _10051_/A vssd1 vssd1 vccd1 vccd1 _11142_/A sky130_fd_sc_hd__or2b_1
XANTENNA__13258__C _14824_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput77 _12013_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[13] sky130_fd_sc_hd__buf_2
X_11072_ _10834_/X _12465_/A _11696_/A _12463_/A vssd1 vssd1 vccd1 vccd1 _11258_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_1_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput88 _12265_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[23] sky130_fd_sc_hd__buf_2
Xoutput99 _11748_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[4] sky130_fd_sc_hd__buf_2
X_10023_ _18838_/Q _19392_/Q _19554_/Q _18806_/Q _09782_/A _09979_/X vssd1 vssd1 vccd1
+ vccd1 _10023_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14900_ _14900_/A _14900_/B vssd1 vssd1 vccd1 vccd1 _14960_/A sky130_fd_sc_hd__and2_1
XANTENNA__09922__C1 _09854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17027__A _17049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_1_clock clkbuf_1_0_1_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_15880_ _16847_/A _17391_/A vssd1 vssd1 vccd1 vccd1 _15937_/A sky130_fd_sc_hd__or2_2
XFILLER_49_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input23_A io_dbus_rdata[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14831_ _14811_/X _14826_/X _14829_/X _14830_/X vssd1 vssd1 vccd1 vccd1 _16673_/A
+ sky130_fd_sc_hd__o31a_4
XFILLER_5_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17461__S _17461_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17550_ _17550_/A vssd1 vssd1 vccd1 vccd1 _19634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14762_ _14761_/X _18590_/Q _14762_/S vssd1 vssd1 vccd1 vccd1 _14763_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11974_ _10461_/A _18502_/Q _12060_/A vssd1 vssd1 vccd1 vccd1 _12011_/A sky130_fd_sc_hd__mux2_8
XANTENNA_clkbuf_leaf_57_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17212__A1 _13334_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16501_ _16134_/X _19210_/Q _16501_/S vssd1 vssd1 vccd1 vccd1 _16502_/A sky130_fd_sc_hd__mux2_1
X_13713_ _13801_/A vssd1 vssd1 vccd1 vccd1 _13796_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10925_ _10973_/A _10925_/B vssd1 vssd1 vccd1 vccd1 _10925_/X sky130_fd_sc_hd__or2_1
X_17481_ _19604_/Q _16664_/X _17485_/S vssd1 vssd1 vccd1 vccd1 _17482_/A sky130_fd_sc_hd__mux2_1
X_14693_ _14587_/A _14648_/X _14680_/X input57/X vssd1 vssd1 vccd1 vccd1 _14694_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19220_ _19541_/CLK _19220_/D vssd1 vssd1 vccd1 vccd1 _19220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16432_ _16488_/A vssd1 vssd1 vccd1 vccd1 _16501_/S sky130_fd_sc_hd__buf_6
X_13644_ _12510_/B _12446_/B _13689_/S vssd1 vssd1 vccd1 vccd1 _13996_/B sky130_fd_sc_hd__mux2_2
XFILLER_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10856_ _09927_/A _10846_/X _10855_/X _09306_/A _18431_/Q vssd1 vssd1 vccd1 vccd1
+ _12466_/A sky130_fd_sc_hd__a32o_4
XANTENNA__12588__A1 _19676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12588__B2 _19486_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19151_ _19700_/CLK _19151_/D vssd1 vssd1 vccd1 vccd1 _19151_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16363_ _19148_/Q _15494_/X _16369_/S vssd1 vssd1 vccd1 vccd1 _16364_/A sky130_fd_sc_hd__mux2_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13682_/S vssd1 vssd1 vccd1 vccd1 _13657_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__09453__A1 _09695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _10895_/A _10787_/B vssd1 vssd1 vccd1 vccd1 _10787_/X sky130_fd_sc_hd__or2_1
X_18102_ _19821_/Q _18102_/B _18102_/C vssd1 vssd1 vccd1 vccd1 _18104_/B sky130_fd_sc_hd__and3_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _18709_/Q _15203_/X _15322_/S vssd1 vssd1 vccd1 vccd1 _15315_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _12526_/A vssd1 vssd1 vccd1 vccd1 _12583_/A sky130_fd_sc_hd__clkbuf_2
X_19082_ _19082_/CLK _19082_/D vssd1 vssd1 vccd1 vccd1 _19082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16294_ _16045_/X _19118_/Q _16296_/S vssd1 vssd1 vccd1 vccd1 _16295_/A sky130_fd_sc_hd__mux2_1
X_18033_ _18033_/A _18033_/B _18033_/C vssd1 vssd1 vccd1 vccd1 _19797_/D sky130_fd_sc_hd__nor3_1
X_15245_ _15264_/S vssd1 vssd1 vccd1 vccd1 _15260_/S sky130_fd_sc_hd__buf_2
X_12457_ _19759_/Q _12186_/X _12454_/X _12456_/X vssd1 vssd1 vccd1 vccd1 _12457_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_output91_A _12333_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ _11423_/A _12537_/B vssd1 vssd1 vccd1 vccd1 _12670_/C sky130_fd_sc_hd__nor2_1
XANTENNA__10446__S0 _11112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15176_ _18662_/Q _15175_/X _15185_/S vssd1 vssd1 vccd1 vccd1 _15177_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12388_ _12388_/A _12410_/B vssd1 vssd1 vccd1 vccd1 _12388_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12353__B _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14127_ _13714_/X _14128_/B _14125_/X _14126_/X vssd1 vssd1 vccd1 vccd1 _14127_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11339_ _11343_/B _11339_/B _11339_/C _13526_/C vssd1 vssd1 vccd1 vccd1 _11339_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_114_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10771__B1 _10797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18935_ _19555_/CLK _18935_/D vssd1 vssd1 vccd1 vccd1 _18935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14058_ _13937_/X _14057_/B _14040_/X vssd1 vssd1 vccd1 vccd1 _14058_/X sky130_fd_sc_hd__o21a_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13009_ _18315_/Q _13004_/C _13008_/Y vssd1 vssd1 vccd1 vccd1 _18315_/D sky130_fd_sc_hd__o21a_1
XANTENNA__10749__S1 _10670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18866_ _19550_/CLK _18866_/D vssd1 vssd1 vccd1 vccd1 _18866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17817_ _17817_/A vssd1 vssd1 vccd1 vccd1 _19710_/D sky130_fd_sc_hd__clkbuf_1
X_18797_ _19223_/CLK _18797_/D vssd1 vssd1 vccd1 vccd1 _18797_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10601__B _10601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17748_ _13376_/X _17747_/Y _17762_/S vssd1 vssd1 vccd1 vccd1 _17748_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17679_ _17683_/A _17683_/C vssd1 vssd1 vccd1 vccd1 _17679_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__17754__A2 _13387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10921__S1 _10920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19418_ _19612_/CLK _19418_/D vssd1 vssd1 vccd1 vccd1 _19418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19349_ _19414_/CLK _19349_/D vssd1 vssd1 vccd1 vccd1 _19349_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10329__A _10329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09102_ _09125_/A vssd1 vssd1 vccd1 vccd1 _11317_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15517__A1 _15516_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10437__S0 _11112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17546__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_132_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _18471_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09935_ _10132_/A vssd1 vssd1 vccd1 vccd1 _09936_/A sky130_fd_sc_hd__buf_2
XFILLER_98_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09866_ _09866_/A vssd1 vssd1 vccd1 vccd1 _09866_/X sky130_fd_sc_hd__buf_4
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13094__B _13104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_147_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19696_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_85_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09797_ _19621_/Q _19459_/Q _18905_/Q _18675_/Q _09976_/A _09763_/A vssd1 vssd1 vccd1
+ vccd1 _09798_/B sky130_fd_sc_hd__mux4_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16686__A _16686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11165__S1 _10306_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09683__A1 _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_clock clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__17745__A2 _13364_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10710_ _10710_/A vssd1 vssd1 vccd1 vccd1 _10711_/A sky130_fd_sc_hd__buf_6
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16953__A0 _16790_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _18572_/Q vssd1 vssd1 vccd1 vccd1 _14557_/A sky130_fd_sc_hd__buf_2
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10641_ _19637_/Q _19054_/Q _19091_/Q _18697_/Q _10631_/X _10634_/X vssd1 vssd1 vccd1
+ vccd1 _10641_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10239__A _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13360_ _18260_/Q _12651_/A _12528_/A _19849_/Q vssd1 vssd1 vccd1 vccd1 _13360_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15508__A1 _15506_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10572_ _10475_/A _10571_/X _09434_/A vssd1 vssd1 vccd1 vccd1 _10572_/X sky130_fd_sc_hd__o21a_1
XFILLER_42_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12311_ _12309_/Y _12311_/B vssd1 vssd1 vccd1 vccd1 _12313_/A sky130_fd_sc_hd__and2b_2
X_13291_ _19838_/Q _12735_/A _12753_/A _19774_/Q vssd1 vssd1 vccd1 vccd1 _13291_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15030_ _14744_/X _15029_/X _14842_/X vssd1 vssd1 vccd1 vccd1 _15030_/X sky130_fd_sc_hd__o21a_1
X_12242_ _12242_/A vssd1 vssd1 vccd1 vccd1 _12244_/B sky130_fd_sc_hd__buf_4
XANTENNA__13269__B _18632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12173_ _12173_/A _12323_/A vssd1 vssd1 vccd1 vccd1 _12173_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09763__A _09763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11124_ _19610_/Q _19448_/Q _18894_/Q _18664_/Q _10279_/S _10245_/X vssd1 vssd1 vccd1
+ vccd1 _11124_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16981_ _16981_/A vssd1 vssd1 vccd1 vccd1 _19397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13285__A _18281_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18720_ _19647_/CLK _18720_/D vssd1 vssd1 vccd1 vccd1 _18720_/Q sky130_fd_sc_hd__dfxtp_1
X_15932_ _15932_/A vssd1 vssd1 vccd1 vccd1 _18967_/D sky130_fd_sc_hd__clkbuf_1
X_11055_ _18753_/Q _18982_/Q _18913_/Q _19211_/Q _10805_/A _10725_/A vssd1 vssd1 vccd1
+ vccd1 _11056_/B sky130_fd_sc_hd__mux4_1
XFILLER_114_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10006_ _10006_/A vssd1 vssd1 vccd1 vccd1 _11269_/A sky130_fd_sc_hd__inv_2
X_15863_ _14996_/X _18937_/Q _15863_/S vssd1 vssd1 vccd1 vccd1 _15864_/A sky130_fd_sc_hd__mux2_1
X_18651_ _19436_/CLK _18651_/D vssd1 vssd1 vccd1 vccd1 _18651_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11517__B _11517_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14247__A1 _14246_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15704__S _15708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14814_ _18435_/Q _14839_/S _14813_/X _14980_/A vssd1 vssd1 vccd1 vccd1 _14814_/X
+ sky130_fd_sc_hd__o211a_1
X_17602_ _17602_/A vssd1 vssd1 vccd1 vccd1 _19658_/D sky130_fd_sc_hd__clkbuf_1
X_15794_ _15009_/X _18906_/Q _15802_/S vssd1 vssd1 vccd1 vccd1 _15795_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18582_ _18585_/CLK _18582_/D vssd1 vssd1 vccd1 vccd1 _18582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17533_ _19628_/Q _16740_/X _17533_/S vssd1 vssd1 vccd1 vccd1 _17534_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14745_ _14743_/A _17621_/A _14744_/X vssd1 vssd1 vccd1 vccd1 _14745_/Y sky130_fd_sc_hd__o21ai_1
X_11957_ _19739_/Q _11957_/B vssd1 vssd1 vccd1 vccd1 _11957_/Y sky130_fd_sc_hd__xnor2_1
X_17464_ _17520_/A vssd1 vssd1 vccd1 vccd1 _17533_/S sky130_fd_sc_hd__buf_6
X_10908_ _09168_/A _10907_/X _10923_/A vssd1 vssd1 vccd1 vccd1 _10908_/X sky130_fd_sc_hd__a21o_1
X_14676_ _14575_/A _14633_/X _14622_/X input51/X vssd1 vssd1 vccd1 vccd1 _14677_/B
+ sky130_fd_sc_hd__a22o_1
X_11888_ _18358_/Q _18357_/Q _11888_/C _11888_/D vssd1 vssd1 vccd1 vccd1 _11962_/D
+ sky130_fd_sc_hd__and4_2
X_19203_ _19427_/CLK _19203_/D vssd1 vssd1 vccd1 vccd1 _19203_/Q sky130_fd_sc_hd__dfxtp_1
X_16415_ _16415_/A vssd1 vssd1 vccd1 vccd1 _16424_/S sky130_fd_sc_hd__clkbuf_8
X_13627_ _13619_/X _13626_/X _13759_/S vssd1 vssd1 vccd1 vccd1 _13627_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17395_ _17395_/A vssd1 vssd1 vccd1 vccd1 _19565_/D sky130_fd_sc_hd__clkbuf_1
X_10839_ _10887_/A _10838_/X _10791_/A vssd1 vssd1 vccd1 vccd1 _10839_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12067__C _19743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09938__A _09969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16346_ _16346_/A vssd1 vssd1 vccd1 vccd1 _19141_/D sky130_fd_sc_hd__clkbuf_1
X_19134_ _19648_/CLK _19134_/D vssd1 vssd1 vccd1 vccd1 _19134_/Q sky130_fd_sc_hd__dfxtp_1
X_13558_ _13558_/A vssd1 vssd1 vccd1 vccd1 _18423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19065_ _19660_/CLK _19065_/D vssd1 vssd1 vccd1 vccd1 _19065_/Q sky130_fd_sc_hd__dfxtp_1
X_12509_ _13742_/S vssd1 vssd1 vccd1 vccd1 _13747_/S sky130_fd_sc_hd__clkbuf_2
X_16277_ _16125_/X _19111_/Q _16279_/S vssd1 vssd1 vccd1 vccd1 _16278_/A sky130_fd_sc_hd__mux2_1
X_13489_ _18403_/Q _12656_/B _13497_/S vssd1 vssd1 vccd1 vccd1 _13490_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18016_ _19790_/Q _18014_/B _18015_/Y vssd1 vssd1 vccd1 vccd1 _19790_/D sky130_fd_sc_hd__o21a_1
X_15228_ _15228_/A vssd1 vssd1 vccd1 vccd1 _18678_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12194__C1 _12193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17366__S _17374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11092__S0 _09449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15159_ _16661_/A vssd1 vssd1 vccd1 vccd1 _15159_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_141_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_64_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19871_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_141_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17890__A _17890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ _09277_/A _09710_/X _09719_/X _09284_/A _18452_/Q vssd1 vssd1 vccd1 vccd1
+ _11222_/A sky130_fd_sc_hd__a32o_4
XANTENNA__11708__A _11749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18918_ _19442_/CLK _18918_/D vssd1 vssd1 vccd1 vccd1 _18918_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10612__A _19693_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09651_ _10309_/A _09651_/B vssd1 vssd1 vccd1 vccd1 _09651_/X sky130_fd_sc_hd__or2_1
X_18849_ _19534_/CLK _18849_/D vssd1 vssd1 vccd1 vccd1 _18849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09582_ _11110_/S vssd1 vssd1 vccd1 vccd1 _09583_/A sky130_fd_sc_hd__buf_4
XFILLER_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_79_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19628_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17188__A0 _18440_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10578__A3 _10577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19550_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_136_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14174__B1 _15123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17276__S _17280_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09583__A _09583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09918_ _18776_/Q _19005_/Q _18936_/Q _19234_/Q _09914_/A _09770_/X vssd1 vssd1 vccd1
+ vccd1 _09919_/B sky130_fd_sc_hd__mux4_1
XANTENNA__11618__A _11618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09849_ _09843_/X _09845_/X _09847_/X _09919_/A _09217_/A vssd1 vssd1 vccd1 vccd1
+ _09854_/B sky130_fd_sc_hd__o221a_1
XFILLER_19_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15524__S _15536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12860_ _12863_/B _12863_/C _12859_/Y vssd1 vssd1 vccd1 vccd1 _18267_/D sky130_fd_sc_hd__o21a_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _11811_/A _13630_/A vssd1 vssd1 vccd1 vccd1 _11811_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17179__A0 _19480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _12791_/A _12791_/B vssd1 vssd1 vccd1 vccd1 _12791_/X sky130_fd_sc_hd__or2_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09656__A1 _09689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _18562_/Q _12763_/X _14529_/Y _14514_/X vssd1 vssd1 vccd1 vccd1 _18530_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _10834_/X _18494_/Q _11840_/A vssd1 vssd1 vccd1 vccd1 _11784_/A sky130_fd_sc_hd__mux2_4
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10671__C1 _10670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _18502_/Q _17878_/A _14465_/S vssd1 vssd1 vccd1 vccd1 _14462_/A sky130_fd_sc_hd__mux2_1
X_11673_ _18343_/Q _18338_/Q vssd1 vssd1 vccd1 vccd1 _11673_/Y sky130_fd_sc_hd__nand2_1
XFILLER_144_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16355__S _16355_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16200_ _16200_/A vssd1 vssd1 vccd1 vccd1 _19072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13412_ _13297_/X _13403_/Y _13411_/X _13306_/X hold3/X vssd1 vssd1 vccd1 vccd1 _13412_/X
+ sky130_fd_sc_hd__a32o_4
X_17180_ _17180_/A vssd1 vssd1 vccd1 vccd1 _19480_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09758__A _10094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ _10750_/A _10624_/B vssd1 vssd1 vccd1 vccd1 _10624_/X sky130_fd_sc_hd__or2_1
XFILLER_139_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14392_ _18476_/Q vssd1 vssd1 vccd1 vccd1 _17701_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16131_ _16841_/A vssd1 vssd1 vccd1 vccd1 _16131_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13343_ _19846_/Q _12736_/A _13340_/X _13342_/X vssd1 vssd1 vccd1 vccd1 _13343_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10555_ _10554_/B _12476_/B vssd1 vssd1 vccd1 vccd1 _10556_/B sky130_fd_sc_hd__and2b_1
X_16062_ _16061_/X _19022_/Q _16065_/S vssd1 vssd1 vccd1 vccd1 _16063_/A sky130_fd_sc_hd__mux2_1
X_13274_ _19869_/Q _12525_/X _12753_/X _19773_/Q vssd1 vssd1 vccd1 vccd1 _14859_/C
+ sky130_fd_sc_hd__a22o_2
XFILLER_143_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ _18597_/Q _19286_/Q _10486_/S vssd1 vssd1 vccd1 vccd1 _10486_/X sky130_fd_sc_hd__mux2_1
X_15013_ input19/X _14924_/X _15000_/X vssd1 vssd1 vccd1 vccd1 _15013_/Y sky130_fd_sc_hd__a21oi_1
X_12225_ _19749_/Q _12002_/X _12224_/Y vssd1 vssd1 vccd1 vccd1 _12225_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12912__A _12997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19821_ _19822_/CLK _19821_/D vssd1 vssd1 vccd1 vccd1 _19821_/Q sky130_fd_sc_hd__dfxtp_1
X_12156_ _14178_/B _12132_/B _12348_/A vssd1 vssd1 vccd1 vccd1 _12157_/B sky130_fd_sc_hd__o21ai_1
XFILLER_151_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14468__A1 _19743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ _11123_/A _11107_/B vssd1 vssd1 vccd1 vccd1 _11107_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19752_ _19755_/CLK _19752_/D vssd1 vssd1 vccd1 vccd1 _19752_/Q sky130_fd_sc_hd__dfxtp_4
X_16964_ _16806_/X _19390_/Q _16964_/S vssd1 vssd1 vccd1 vccd1 _16965_/A sky130_fd_sc_hd__mux2_1
X_12087_ _12036_/A _12064_/A _12064_/B vssd1 vssd1 vccd1 vccd1 _12087_/X sky130_fd_sc_hd__o21ba_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18703_ _19579_/CLK _18703_/D vssd1 vssd1 vccd1 vccd1 _18703_/Q sky130_fd_sc_hd__dfxtp_1
X_15915_ _15937_/A vssd1 vssd1 vccd1 vccd1 _15924_/S sky130_fd_sc_hd__buf_4
X_11038_ _19629_/Q _19046_/Q _19083_/Q _18689_/Q _10663_/A _10364_/A vssd1 vssd1 vccd1
+ vccd1 _11038_/X sky130_fd_sc_hd__mux4_2
X_19683_ _19686_/CLK _19683_/D vssd1 vssd1 vccd1 vccd1 _19683_/Q sky130_fd_sc_hd__dfxtp_2
X_16895_ _16895_/A vssd1 vssd1 vccd1 vccd1 _19359_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18634_ _19081_/CLK _18634_/D vssd1 vssd1 vccd1 vccd1 _18634_/Q sky130_fd_sc_hd__dfxtp_2
X_15846_ _14908_/X _18929_/Q _15852_/S vssd1 vssd1 vccd1 vccd1 _15847_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18565_ _18585_/CLK _18565_/D vssd1 vssd1 vccd1 vccd1 _18565_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_18_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09647__A1 _09562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ _12993_/A _12993_/C _12922_/X vssd1 vssd1 vccd1 vccd1 _12989_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15777_ _15777_/A vssd1 vssd1 vccd1 vccd1 _18898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17516_ _19620_/Q _16715_/X _17518_/S vssd1 vssd1 vccd1 vccd1 _17517_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09742__S1 _10186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14728_ _16645_/A vssd1 vssd1 vccd1 vccd1 _16749_/A sky130_fd_sc_hd__clkbuf_2
X_18496_ _19693_/CLK _18496_/D vssd1 vssd1 vccd1 vccd1 _18496_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17447_ _17447_/A vssd1 vssd1 vccd1 vccd1 _19589_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14659_ _14659_/A vssd1 vssd1 vccd1 vccd1 _18572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11206__A1 _11203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17378_ _17378_/A vssd1 vssd1 vccd1 vccd1 _19558_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12954__A1 _18295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19117_ _19633_/CLK _19117_/D vssd1 vssd1 vccd1 vccd1 _19117_/Q sky130_fd_sc_hd__dfxtp_1
X_16329_ _16096_/X _19134_/Q _16329_/S vssd1 vssd1 vccd1 vccd1 _16330_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19048_ _19633_/CLK _19048_/D vssd1 vssd1 vccd1 vccd1 _19048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_179_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12706__B2 _19480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10193__A1 _09404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14459__A1 _19739_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15120__A2 _15116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13131__A1 _19856_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09703_ _10103_/A _09699_/X _09702_/X vssd1 vssd1 vccd1 vccd1 _09703_/X sky130_fd_sc_hd__a21o_1
XFILLER_114_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13653__A _13653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ _09634_/A vssd1 vssd1 vccd1 vccd1 _09635_/A sky130_fd_sc_hd__buf_2
XFILLER_95_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11693__A1 _18564_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12890__B1 _12869_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09565_ _19530_/Q _19144_/Q _19594_/Q _18750_/Q _09553_/X _09144_/A vssd1 vssd1 vccd1
+ vccd1 _09566_/B sky130_fd_sc_hd__mux4_1
XFILLER_167_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13434__A2 _12665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09496_ _10934_/S vssd1 vssd1 vccd1 vccd1 _10631_/A sky130_fd_sc_hd__buf_4
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16175__S _16183_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11901__A _11901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17333__A0 _16761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11112__S _11112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10340_ _19612_/Q _19450_/Q _18896_/Q _18666_/Q _10129_/S _09723_/A vssd1 vssd1 vccd1
+ vccd1 _10341_/B sky130_fd_sc_hd__mux4_1
XFILLER_164_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10271_ _18833_/Q _19387_/Q _19549_/Q _18801_/Q _11156_/S _09145_/A vssd1 vssd1 vccd1
+ vccd1 _10271_/X sky130_fd_sc_hd__mux4_2
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13370__A1 _19685_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ _12010_/A _13595_/A vssd1 vssd1 vccd1 vccd1 _12013_/A sky130_fd_sc_hd__xor2_4
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17636__A1 _17634_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13961_ _11787_/Y _14070_/A _13951_/X _13960_/Y vssd1 vssd1 vccd1 vccd1 _13961_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14870__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12912_ _12997_/A _12919_/C vssd1 vssd1 vccd1 vccd1 _12912_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15700_ _18864_/Q _15538_/X _15708_/S vssd1 vssd1 vccd1 vccd1 _15701_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13563__A _13563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16680_ _16680_/A vssd1 vssd1 vccd1 vccd1 _16680_/X sky130_fd_sc_hd__buf_2
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13892_ _13883_/X _13890_/X _13970_/S vssd1 vssd1 vccd1 vccd1 _13892_/X sky130_fd_sc_hd__mux2_2
XFILLER_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12843_ _12854_/D vssd1 vssd1 vccd1 vccd1 _12850_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15631_ _15631_/A vssd1 vssd1 vccd1 vccd1 _18833_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13425__A2 _13423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_opt_4_0_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18350_ _18357_/CLK _18350_/D vssd1 vssd1 vccd1 vccd1 _18350_/Q sky130_fd_sc_hd__dfxtp_1
X_15562_ _18807_/Q _15561_/X _15568_/S vssd1 vssd1 vccd1 vccd1 _15563_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _18327_/Q _13130_/A _12735_/A _19848_/Q vssd1 vssd1 vccd1 vccd1 _12774_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09724__S1 _09723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _17301_/A vssd1 vssd1 vccd1 vccd1 _19524_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_6_0_clock clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
X_14513_ _14513_/A _14519_/B vssd1 vssd1 vccd1 vccd1 _14513_/X sky130_fd_sc_hd__or2_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _18353_/Q _11759_/B vssd1 vssd1 vccd1 vccd1 _11726_/B sky130_fd_sc_hd__xor2_1
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18281_ _18402_/CLK _18281_/D vssd1 vssd1 vccd1 vccd1 _18281_/Q sky130_fd_sc_hd__dfxtp_1
X_15493_ _15493_/A vssd1 vssd1 vccd1 vccd1 _18785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16085__S _16097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12907__A _18281_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17232_ _18453_/Q _13387_/X _17235_/S vssd1 vssd1 vccd1 vccd1 _17232_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09488__A _10724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14444_ _14444_/A vssd1 vssd1 vccd1 vccd1 _18494_/D sky130_fd_sc_hd__clkbuf_1
X_11656_ input66/X _12715_/A vssd1 vssd1 vccd1 vccd1 _11999_/A sky130_fd_sc_hd__and2_1
XFILLER_156_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12936__A1 _18289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17163_ _17163_/A vssd1 vssd1 vccd1 vccd1 _19475_/D sky130_fd_sc_hd__clkbuf_1
X_10607_ _09538_/A _10604_/X _10606_/X vssd1 vssd1 vccd1 vccd1 _10607_/X sky130_fd_sc_hd__a21o_1
XFILLER_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17324__A0 _16749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14375_ _18470_/Q vssd1 vssd1 vccd1 vccd1 _14861_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11587_ _11587_/A _11587_/B _11587_/C vssd1 vssd1 vccd1 vccd1 _11831_/A sky130_fd_sc_hd__or3_4
XANTENNA__09801__B2 _18450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16114_ _16114_/A vssd1 vssd1 vccd1 vccd1 _19038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13326_ _18288_/Q _13326_/B vssd1 vssd1 vccd1 vccd1 _13326_/X sky130_fd_sc_hd__and2_1
XFILLER_156_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10538_ _19253_/Q _19024_/Q _18955_/Q _19349_/Q _10604_/S _10367_/A vssd1 vssd1 vccd1
+ vccd1 _10539_/B sky130_fd_sc_hd__mux4_1
X_17094_ _17094_/A vssd1 vssd1 vccd1 vccd1 _19447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16045_ _16755_/A vssd1 vssd1 vccd1 vccd1 _16045_/X sky130_fd_sc_hd__clkbuf_1
X_13257_ _19834_/Q _12736_/X _13256_/X vssd1 vssd1 vccd1 vccd1 _14824_/D sky130_fd_sc_hd__a21o_1
XFILLER_170_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10469_ _19414_/Q _19190_/Q _19707_/Q _19158_/Q _09447_/A _09635_/A vssd1 vssd1 vccd1
+ vccd1 _10469_/X sky130_fd_sc_hd__mux4_1
X_12208_ _12209_/A _14216_/B vssd1 vssd1 vccd1 vccd1 _12210_/A sky130_fd_sc_hd__nor2_1
XFILLER_97_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13188_ _19765_/Q vssd1 vssd1 vccd1 vccd1 _17944_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_124_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19804_ _19804_/CLK _19804_/D vssd1 vssd1 vccd1 vccd1 _19804_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15953__A _17892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _12086_/A _12112_/A _12112_/B vssd1 vssd1 vccd1 vccd1 _12139_/X sky130_fd_sc_hd__o21ba_1
XFILLER_69_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17996_ _19783_/Q _17997_/C _19784_/Q vssd1 vssd1 vccd1 vccd1 _17998_/B sky130_fd_sc_hd__a21oi_1
XFILLER_85_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13113__A1 _17149_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09951__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19735_ _19738_/CLK _19735_/D vssd1 vssd1 vccd1 vccd1 _19735_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16947_ _16781_/X _19382_/Q _16953_/S vssd1 vssd1 vccd1 vccd1 _16948_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19666_ _19786_/CLK _19666_/D vssd1 vssd1 vccd1 vccd1 _19666_/Q sky130_fd_sc_hd__dfxtp_4
X_16878_ _19352_/Q _16683_/X _16880_/S vssd1 vssd1 vccd1 vccd1 _16879_/A sky130_fd_sc_hd__mux2_1
X_18617_ _19628_/CLK _18617_/D vssd1 vssd1 vccd1 vccd1 _18617_/Q sky130_fd_sc_hd__dfxtp_1
X_15829_ _15829_/A vssd1 vssd1 vccd1 vccd1 _18921_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19597_ _19597_/CLK _19597_/D vssd1 vssd1 vccd1 vccd1 _19597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16784__A _16784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09350_ _18978_/Q vssd1 vssd1 vccd1 vccd1 _10712_/A sky130_fd_sc_hd__buf_2
X_18548_ _18548_/CLK _18548_/D vssd1 vssd1 vccd1 vccd1 _18548_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09715__S1 _10080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09281_ _09281_/A vssd1 vssd1 vccd1 vccd1 _09282_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10051__B_N _12491_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18479_ _18510_/CLK _18479_/D vssd1 vssd1 vccd1 vccd1 _18479_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12817__A _18173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09398__A _10944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17819__S _17827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16723__S _16735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10337__A _11185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11168__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10261__S1 _09144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09861__A _09861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11115__B1 _09529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09617_ _11178_/A _09615_/X _09616_/X vssd1 vssd1 vccd1 vccd1 _09617_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15802__S _15802_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10011__S _10011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ _09978_/A _09545_/X _09547_/X vssd1 vssd1 vccd1 vccd1 _09548_/X sky130_fd_sc_hd__a21o_1
XFILLER_169_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09706__S1 _09704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09479_ _10725_/A vssd1 vssd1 vccd1 vccd1 _09480_/A sky130_fd_sc_hd__buf_2
XFILLER_24_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11510_ _13523_/B _14568_/A vssd1 vssd1 vccd1 vccd1 _11628_/A sky130_fd_sc_hd__or2_1
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12490_ _12490_/A vssd1 vssd1 vccd1 vccd1 _12490_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12446__B _12446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11441_ _18415_/Q _18427_/Q vssd1 vssd1 vccd1 vccd1 _11723_/B sky130_fd_sc_hd__nand2_1
XFILLER_138_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14160_ _12096_/B _14070_/A _14158_/X _14159_/Y vssd1 vssd1 vccd1 vccd1 _14160_/X
+ sky130_fd_sc_hd__a22o_1
X_11372_ _11372_/A _11372_/B vssd1 vssd1 vccd1 vccd1 _11479_/A sky130_fd_sc_hd__and2_1
XFILLER_164_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13111_ _18348_/Q _13109_/X _13110_/X _13102_/X vssd1 vssd1 vccd1 vccd1 _18348_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18133__B _19830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11072__A1_N _10834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10323_ _09276_/A _10311_/X _10322_/X _09283_/A _18441_/Q vssd1 vssd1 vccd1 vccd1
+ _11135_/A sky130_fd_sc_hd__a32o_4
X_14091_ _14089_/B _14093_/A vssd1 vssd1 vccd1 vccd1 _14092_/B sky130_fd_sc_hd__and2b_1
XFILLER_106_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12462__A _12462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09547__B1 _09184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input53_A io_ibus_inst[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ _13042_/A vssd1 vssd1 vccd1 vccd1 _18085_/A sky130_fd_sc_hd__buf_2
XFILLER_124_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10254_ _19259_/Q _19030_/Q _18961_/Q _19355_/Q _09794_/A _09697_/A vssd1 vssd1 vccd1
+ vccd1 _10255_/B sky130_fd_sc_hd__mux4_1
XFILLER_133_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17850_ _17850_/A vssd1 vssd1 vccd1 vccd1 _19725_/D sky130_fd_sc_hd__clkbuf_1
X_10185_ _18604_/Q _19293_/Q _10185_/S vssd1 vssd1 vccd1 vccd1 _10186_/B sky130_fd_sc_hd__mux2_1
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16801_ _16800_/X _19324_/Q _16807_/S vssd1 vssd1 vccd1 vccd1 _16802_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17781_ _17781_/A _17781_/B vssd1 vssd1 vccd1 vccd1 _17782_/A sky130_fd_sc_hd__and2_2
XFILLER_93_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14993_ _14990_/Y _14991_/X _14992_/X _14838_/A _14999_/A vssd1 vssd1 vccd1 vccd1
+ _14994_/B sky130_fd_sc_hd__a221o_1
XANTENNA__13293__A _18633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19520_ _19648_/CLK _19520_/D vssd1 vssd1 vccd1 vccd1 _19520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16732_ _19303_/Q _16731_/X _16735_/S vssd1 vssd1 vccd1 vccd1 _16733_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09945__S1 _09881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13944_ _13939_/B _13936_/B _13941_/X _13943_/Y vssd1 vssd1 vccd1 vccd1 _13944_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_127_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19451_ _19452_/CLK _19451_/D vssd1 vssd1 vccd1 vccd1 _19451_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11525__B _12466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16663_ _16663_/A vssd1 vssd1 vccd1 vccd1 _19281_/D sky130_fd_sc_hd__clkbuf_1
X_13875_ _13872_/X _13874_/Y _18428_/Q _13736_/X vssd1 vssd1 vccd1 vccd1 _18428_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18402_ _18402_/CLK _18402_/D vssd1 vssd1 vccd1 vccd1 _18402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12826_ _18257_/Q _12822_/C _12825_/Y vssd1 vssd1 vccd1 vccd1 _18257_/D sky130_fd_sc_hd__o21a_1
X_15614_ _18826_/Q _15519_/X _15614_/S vssd1 vssd1 vccd1 vccd1 _15615_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19382_ _19608_/CLK _19382_/D vssd1 vssd1 vccd1 vccd1 _19382_/Q sky130_fd_sc_hd__dfxtp_1
X_16594_ _16594_/A vssd1 vssd1 vccd1 vccd1 _19252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18333_ _19866_/CLK _18333_/D vssd1 vssd1 vccd1 vccd1 _18333_/Q sky130_fd_sc_hd__dfxtp_1
X_12757_ _12556_/X _12733_/Y _12756_/X _12712_/X _18642_/Q vssd1 vssd1 vccd1 vccd1
+ _12757_/X sky130_fd_sc_hd__a32o_4
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15545_ _16800_/A vssd1 vssd1 vccd1 vccd1 _15545_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16109__A _16819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11749_/A vssd1 vssd1 vccd1 vccd1 _12389_/S sky130_fd_sc_hd__buf_2
X_18264_ _19779_/CLK _18264_/D vssd1 vssd1 vccd1 vccd1 _18264_/Q sky130_fd_sc_hd__dfxtp_1
X_15476_ _15476_/A vssd1 vssd1 vccd1 vccd1 _18779_/D sky130_fd_sc_hd__clkbuf_1
X_12688_ _14582_/A _12734_/A _12688_/C vssd1 vssd1 vccd1 vccd1 _16211_/B sky130_fd_sc_hd__or3_2
XFILLER_30_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15020__A1 _14711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12909__A1 _18281_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17215_ _18448_/Q _13346_/X _17218_/S vssd1 vssd1 vccd1 vccd1 _17215_/X sky130_fd_sc_hd__mux2_1
X_14427_ _18488_/Q _18520_/Q _15087_/S vssd1 vssd1 vccd1 vccd1 _14428_/A sky130_fd_sc_hd__mux2_1
X_11639_ _11639_/A _13583_/B vssd1 vssd1 vccd1 vccd1 _13584_/B sky130_fd_sc_hd__nor2_1
X_18195_ _19852_/Q _18196_/C _18194_/Y vssd1 vssd1 vccd1 vccd1 _19852_/D sky130_fd_sc_hd__o21a_1
XFILLER_128_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16543__S _16547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17146_ _18428_/Q _15258_/X _15255_/B vssd1 vssd1 vccd1 vccd1 _17146_/X sky130_fd_sc_hd__a21o_1
X_14358_ _18464_/Q vssd1 vssd1 vccd1 vccd1 _14786_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13309_ _18365_/Q _13319_/B vssd1 vssd1 vccd1 vccd1 _13309_/X sky130_fd_sc_hd__or2_1
XFILLER_155_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17077_ _17134_/S vssd1 vssd1 vccd1 vccd1 _17086_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_171_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14289_ _14289_/A _14289_/B vssd1 vssd1 vccd1 vccd1 _14289_/X sky130_fd_sc_hd__or2_1
XANTENNA__12372__A _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10491__S1 _10238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13187__B _18624_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16028_ _16028_/A vssd1 vssd1 vccd1 vccd1 _19011_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17374__S _17374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09681__A _09681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17979_ _19778_/Q _19777_/Q _17979_/C vssd1 vssd1 vccd1 vccd1 _17981_/B sky130_fd_sc_hd__and3_1
X_19718_ _19718_/CLK _19718_/D vssd1 vssd1 vccd1 vccd1 _19718_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11716__A _11716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19649_ _19810_/CLK _19649_/D vssd1 vssd1 vccd1 vccd1 _19649_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11435__B _12555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09402_ _09402_/A vssd1 vssd1 vccd1 vccd1 _09403_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09333_ _09969_/A vssd1 vssd1 vccd1 vccd1 _09819_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_34_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11451__A _11716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09264_ _18529_/Q vssd1 vssd1 vccd1 vccd1 _16138_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_138_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09195_ _10875_/A vssd1 vssd1 vccd1 vccd1 _10622_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09856__A _09856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12282__A _12282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16689__A _16689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09591__A _10242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11990_ _19671_/Q _11989_/X _11790_/X vssd1 vssd1 vccd1 vccd1 _11990_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10941_ _18756_/Q _18985_/Q _18916_/Q _19214_/Q _09336_/A _10940_/X vssd1 vssd1 vccd1
+ vccd1 _10942_/B sky130_fd_sc_hd__mux4_2
XFILLER_17_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10311__A1 _09214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13660_ _13657_/X _13659_/X _13775_/S vssd1 vssd1 vccd1 vccd1 _13833_/B sky130_fd_sc_hd__mux2_1
X_10872_ _19602_/Q _19440_/Q _18886_/Q _18656_/Q _10664_/S _10365_/A vssd1 vssd1 vccd1
+ vccd1 _10873_/B sky130_fd_sc_hd__mux4_1
XFILLER_72_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12611_ _12930_/C _13404_/B _12609_/X _12610_/X vssd1 vssd1 vccd1 vccd1 _12611_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _13657_/S vssd1 vssd1 vccd1 vccd1 _13724_/B sky130_fd_sc_hd__buf_2
XFILLER_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _15330_/A vssd1 vssd1 vccd1 vccd1 _18716_/D sky130_fd_sc_hd__clkbuf_1
X_12542_ _19675_/Q _12624_/A _13222_/S _19485_/Q vssd1 vssd1 vccd1 vccd1 _12542_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15261_ _15261_/A vssd1 vssd1 vccd1 vccd1 _18687_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17459__S _17461_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12473_ _12473_/A _12483_/B vssd1 vssd1 vccd1 vccd1 _12473_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__16363__S _16369_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14212_ _14212_/A _14216_/A vssd1 vssd1 vccd1 vccd1 _14212_/Y sky130_fd_sc_hd__nand2_1
X_17000_ _17000_/A vssd1 vssd1 vccd1 vccd1 _19405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11424_ _11821_/A _12530_/A _12686_/A _12537_/B vssd1 vssd1 vccd1 vccd1 _12532_/A
+ sky130_fd_sc_hd__nor4_1
XFILLER_126_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15192_ _18667_/Q _15191_/X _15201_/S vssd1 vssd1 vccd1 vccd1 _15193_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14143_ _14140_/B _14138_/B _13862_/A _14141_/X _14142_/X vssd1 vssd1 vccd1 vccd1
+ _14143_/X sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_53_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11355_ _11362_/A vssd1 vssd1 vccd1 vccd1 _11355_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12192__A _19679_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10306_ _10306_/A vssd1 vssd1 vccd1 vccd1 _10306_/X sky130_fd_sc_hd__clkbuf_4
X_18951_ _19702_/CLK _18951_/D vssd1 vssd1 vccd1 vccd1 _18951_/Q sky130_fd_sc_hd__dfxtp_1
X_14074_ _14075_/B _14074_/B vssd1 vssd1 vccd1 vccd1 _14078_/B sky130_fd_sc_hd__nand2_1
XFILLER_140_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11286_ _11205_/Y _11284_/C _13585_/A vssd1 vssd1 vccd1 vccd1 _11286_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__09615__S0 _09729_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17902_ _19752_/Q vssd1 vssd1 vccd1 vccd1 _17902_/Y sky130_fd_sc_hd__inv_2
X_13025_ _13034_/A _13025_/B _13025_/C vssd1 vssd1 vccd1 vccd1 _18320_/D sky130_fd_sc_hd__nor3_1
XFILLER_117_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10237_ _10651_/A vssd1 vssd1 vccd1 vccd1 _10238_/A sky130_fd_sc_hd__clkbuf_4
X_18882_ _19699_/CLK _18882_/D vssd1 vssd1 vccd1 vccd1 _18882_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10225__S1 _09486_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17833_ _17833_/A vssd1 vssd1 vccd1 vccd1 _19717_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10168_ _18835_/Q _19389_/Q _19551_/Q _18803_/Q _10076_/S _09979_/A vssd1 vssd1 vccd1
+ vccd1 _10168_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15008__A _16721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17764_ _17764_/A vssd1 vssd1 vccd1 vccd1 _19688_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10440__A _10447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14976_ _14975_/X _18608_/Q _14997_/S vssd1 vssd1 vccd1 vccd1 _14977_/A sky130_fd_sc_hd__mux2_1
X_10099_ _12489_/C _10098_/X vssd1 vssd1 vccd1 vccd1 _10100_/A sky130_fd_sc_hd__or2b_1
XFILLER_19_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19503_ _19631_/CLK _19503_/D vssd1 vssd1 vccd1 vccd1 _19503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16715_ _16715_/A vssd1 vssd1 vccd1 vccd1 _16715_/X sky130_fd_sc_hd__buf_2
X_13927_ _13927_/A vssd1 vssd1 vccd1 vccd1 _13927_/X sky130_fd_sc_hd__clkbuf_2
X_17695_ _19675_/Q _17694_/X _17718_/S vssd1 vssd1 vccd1 vccd1 _17696_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17766__B1 _18488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15442__S _15448_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19434_ _19727_/CLK _19434_/D vssd1 vssd1 vccd1 vccd1 _19434_/Q sky130_fd_sc_hd__dfxtp_1
X_16646_ _19276_/Q _16645_/X _16655_/S vssd1 vssd1 vccd1 vccd1 _16647_/A sky130_fd_sc_hd__mux2_1
X_13858_ _14320_/A _13913_/S vssd1 vssd1 vccd1 vccd1 _13858_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12809_ _12851_/A _12809_/B _12809_/C vssd1 vssd1 vccd1 vccd1 _18253_/D sky130_fd_sc_hd__nor3_1
X_19365_ _19591_/CLK _19365_/D vssd1 vssd1 vccd1 vccd1 _19365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12367__A _13388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16577_ _19244_/Q vssd1 vssd1 vccd1 vccd1 _16578_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_37_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13789_ _13789_/A vssd1 vssd1 vccd1 vccd1 _13879_/S sky130_fd_sc_hd__buf_2
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10066__B1 _09892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18316_ _18330_/CLK _18316_/D vssd1 vssd1 vccd1 vccd1 _18316_/Q sky130_fd_sc_hd__dfxtp_1
X_15528_ _15528_/A vssd1 vssd1 vccd1 vccd1 _18796_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19296_ _19329_/CLK _19296_/D vssd1 vssd1 vccd1 vccd1 _19296_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_3_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__09471__A2 _09461_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18247_ _19871_/Q _18247_/B _18247_/C vssd1 vssd1 vccd1 vccd1 _18249_/B sky130_fd_sc_hd__and3_1
XANTENNA__16273__S _16279_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15459_ _18772_/Q _15200_/X _15459_/S vssd1 vssd1 vccd1 vccd1 _15460_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09676__A _09735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18178_ _18197_/A _18183_/C vssd1 vssd1 vccd1 vccd1 _18178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17129_ _17129_/A vssd1 vssd1 vccd1 vccd1 _19463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13307__B2 _18634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ _09951_/A _12495_/C vssd1 vssd1 vccd1 vccd1 _11225_/B sky130_fd_sc_hd__or2b_1
XFILLER_131_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18246__A1 _18247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15617__S _15625_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09882_ _19428_/Q _19204_/Q _19721_/Q _19172_/Q _09809_/X _09881_/X vssd1 vssd1 vccd1
+ vccd1 _09882_/X sky130_fd_sc_hd__mux4_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17832__S _17838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12277__A _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ _09621_/A vssd1 vssd1 vccd1 vccd1 _09317_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18182__B1 _19848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09289__C _18575_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09247_ _09247_/A vssd1 vssd1 vccd1 vccd1 _09248_/A sky130_fd_sc_hd__buf_4
XANTENNA__16183__S _16183_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09586__A _10331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09178_ _10996_/A vssd1 vssd1 vccd1 vccd1 _09179_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16911__S _16913_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11140_ _11230_/A _11234_/A _11230_/C _10197_/A _11139_/X vssd1 vssd1 vccd1 vccd1
+ _11227_/C sky130_fd_sc_hd__a311o_1
Xclkbuf_4_5_0_clock clkbuf_4_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_116_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15527__S _15536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput78 _12041_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[14] sky130_fd_sc_hd__buf_2
X_11071_ _11024_/X _11257_/A _11254_/A vssd1 vssd1 vccd1 vccd1 _11071_/X sky130_fd_sc_hd__a21o_1
XFILLER_131_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput89 _12290_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[24] sky130_fd_sc_hd__buf_2
XFILLER_89_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10022_ _10022_/A _10022_/B vssd1 vssd1 vccd1 vccd1 _10022_/X sky130_fd_sc_hd__or2_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14830_ input2/X _14801_/A _14804_/A vssd1 vssd1 vccd1 vccd1 _14830_/X sky130_fd_sc_hd__a21o_1
XFILLER_64_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11075__B _12468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input16_A io_dbus_rdata[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17748__A0 _13376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14761_ _16758_/A vssd1 vssd1 vccd1 vccd1 _14761_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11973_ _14089_/B _11973_/B vssd1 vssd1 vccd1 vccd1 _11975_/A sky130_fd_sc_hd__xnor2_4
XFILLER_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16500_ _16500_/A vssd1 vssd1 vccd1 vccd1 _19209_/D sky130_fd_sc_hd__clkbuf_1
X_10924_ _19631_/Q _19048_/Q _19085_/Q _18691_/Q _10919_/X _10920_/X vssd1 vssd1 vccd1
+ vccd1 _10925_/B sky130_fd_sc_hd__mux4_2
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13712_ _13712_/A _13712_/B _13720_/B vssd1 vssd1 vccd1 vccd1 _13801_/A sky130_fd_sc_hd__or3b_1
XFILLER_72_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17480_ _17480_/A vssd1 vssd1 vccd1 vccd1 _19603_/D sky130_fd_sc_hd__clkbuf_1
X_14692_ _14692_/A vssd1 vssd1 vccd1 vccd1 _18583_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16431_ _16920_/B _17783_/B vssd1 vssd1 vccd1 vccd1 _16488_/A sky130_fd_sc_hd__nand2_4
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13643_ _13643_/A vssd1 vssd1 vccd1 vccd1 _13689_/S sky130_fd_sc_hd__clkbuf_2
X_10855_ _09409_/A _10848_/X _10850_/X _10854_/X _09391_/A vssd1 vssd1 vccd1 vccd1
+ _10855_/X sky130_fd_sc_hd__a311o_2
XANTENNA__12037__B2 _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12187__A _19747_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16882__A _16904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09989__B1 _09988_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19150_ _19699_/CLK _19150_/D vssd1 vssd1 vccd1 vccd1 _19150_/Q sky130_fd_sc_hd__dfxtp_1
X_16362_ _16362_/A vssd1 vssd1 vccd1 vccd1 _19147_/D sky130_fd_sc_hd__clkbuf_1
X_13574_ _13643_/A vssd1 vssd1 vccd1 vccd1 _13682_/S sky130_fd_sc_hd__buf_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11796__A0 _19664_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10786_ _19247_/Q _19018_/Q _18949_/Q _19343_/Q _10711_/A _10785_/X vssd1 vssd1 vccd1
+ vccd1 _10787_/B sky130_fd_sc_hd__mux4_2
XFILLER_12_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18101_ _18102_/B _18102_/C _18100_/Y vssd1 vssd1 vccd1 vccd1 _19820_/D sky130_fd_sc_hd__o21a_1
XFILLER_40_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10599__B2 _18435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12525_ _12651_/A vssd1 vssd1 vccd1 vccd1 _12525_/X sky130_fd_sc_hd__clkbuf_2
X_15313_ _15324_/A vssd1 vssd1 vccd1 vccd1 _15322_/S sky130_fd_sc_hd__buf_4
X_16293_ _16293_/A vssd1 vssd1 vccd1 vccd1 _19117_/D sky130_fd_sc_hd__clkbuf_1
X_19081_ _19081_/CLK _19081_/D vssd1 vssd1 vccd1 vccd1 _19081_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18032_ _18031_/B _18031_/C _19797_/Q vssd1 vssd1 vccd1 vccd1 _18033_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__09496__A _10934_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12456_ _12196_/X _12455_/Y _11997_/X vssd1 vssd1 vccd1 vccd1 _12456_/X sky130_fd_sc_hd__a21o_1
X_15244_ _12671_/X _15241_/X _15243_/Y vssd1 vssd1 vccd1 vccd1 _15264_/S sky130_fd_sc_hd__o21a_1
XFILLER_173_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12634__B _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11407_ _18549_/Q _18547_/Q _18546_/Q _18548_/Q vssd1 vssd1 vccd1 vccd1 _12537_/B
+ sky130_fd_sc_hd__or4b_2
X_15175_ _16677_/A vssd1 vssd1 vccd1 vccd1 _15175_/X sky130_fd_sc_hd__clkbuf_2
X_12387_ _19755_/Q _19756_/Q _12387_/C vssd1 vssd1 vccd1 vccd1 _12410_/B sky130_fd_sc_hd__and3_1
XFILLER_126_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output84_A _11624_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14126_ _14126_/A _14126_/B vssd1 vssd1 vccd1 vccd1 _14126_/X sky130_fd_sc_hd__or2_1
X_11338_ _11338_/A vssd1 vssd1 vccd1 vccd1 _13526_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_98_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10771__A1 _10634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18934_ _19003_/CLK _18934_/D vssd1 vssd1 vccd1 vccd1 _18934_/Q sky130_fd_sc_hd__dfxtp_1
X_14057_ _14059_/B _14057_/B vssd1 vssd1 vccd1 vccd1 _14062_/B sky130_fd_sc_hd__and2_1
X_11269_ _11269_/A _11269_/B _11269_/C vssd1 vssd1 vccd1 vccd1 _11271_/A sky130_fd_sc_hd__nand3_1
XFILLER_95_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13008_ _13049_/A _13015_/C vssd1 vssd1 vccd1 vccd1 _13008_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18865_ _19581_/CLK _18865_/D vssd1 vssd1 vccd1 vccd1 _18865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15961__A _16503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17816_ _15184_/X _19710_/Q _17816_/S vssd1 vssd1 vccd1 vccd1 _17817_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18796_ _19608_/CLK _18796_/D vssd1 vssd1 vccd1 vccd1 _18796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12276__A1 _19751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17747_ _17751_/A _17751_/C vssd1 vssd1 vccd1 vccd1 _17747_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__16268__S _16268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14959_ _18447_/Q _15018_/A _14958_/X _14980_/A vssd1 vssd1 vccd1 vccd1 _14959_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_35_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17678_ _17678_/A vssd1 vssd1 vccd1 vccd1 _19672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19417_ _19710_/CLK _19417_/D vssd1 vssd1 vccd1 vccd1 _19417_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17888__A _17890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16629_ _19270_/Q vssd1 vssd1 vccd1 vccd1 _16630_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15900__S _15902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19348_ _19659_/CLK _19348_/D vssd1 vssd1 vccd1 vccd1 _19348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09101_ _11534_/B _14519_/A _11468_/B vssd1 vssd1 vccd1 vccd1 _11495_/B sky130_fd_sc_hd__or3_2
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19279_ _19601_/CLK _19279_/D vssd1 vssd1 vccd1 vccd1 _19279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14725__A0 _11022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17827__S _17827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10345__A _18441_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15347__S _15351_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09934_ _19426_/Q _19202_/Q _19719_/Q _19170_/Q _09866_/X _09869_/X vssd1 vssd1 vccd1
+ vccd1 _09934_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12560__A input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ _09865_/A vssd1 vssd1 vccd1 vccd1 _09866_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__13375__B _15018_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input8_A io_dbus_rdata[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11176__A _11185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17562__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10080__A _10080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _10153_/S vssd1 vssd1 vccd1 vccd1 _09976_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15453__A1 _15191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11904__A _19668_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10640_ _10640_/A _10640_/B vssd1 vssd1 vccd1 vccd1 _10640_/Y sky130_fd_sc_hd__nor2_1
XFILLER_167_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18155__B1 _19839_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10571_ _19638_/Q _19055_/Q _19092_/Q _18698_/Q _11088_/S _10559_/A vssd1 vssd1 vccd1
+ vccd1 _10571_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12735__A _12735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12310_ _12310_/A _12310_/B vssd1 vssd1 vccd1 vccd1 _12311_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13290_ _18317_/Q _12663_/X _12651_/X _18247_/B vssd1 vssd1 vccd1 vccd1 _14873_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09818__S0 _09803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12241_ _12241_/A _12241_/B vssd1 vssd1 vccd1 vccd1 _12242_/A sky130_fd_sc_hd__and2_1
XANTENNA__14950__A _16705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12172_ _13524_/B _12277_/B vssd1 vssd1 vccd1 vccd1 _12172_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11123_ _11123_/A _11123_/B vssd1 vssd1 vccd1 vccd1 _11123_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13566__A _15116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17038__A _17049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16980_ _16829_/X _19397_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16981_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15931_ _14975_/X _18967_/Q _15935_/S vssd1 vssd1 vccd1 vccd1 _15932_/A sky130_fd_sc_hd__mux2_1
X_11054_ _19403_/Q _19179_/Q _19696_/Q _19147_/Q _10932_/S _10772_/A vssd1 vssd1 vccd1
+ vccd1 _11054_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10505__A1 _09412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17472__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11086__A _11097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ _11272_/A _10005_/B vssd1 vssd1 vccd1 vccd1 _10006_/A sky130_fd_sc_hd__or2_1
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18650_ _19081_/CLK _18650_/D vssd1 vssd1 vccd1 vccd1 _18650_/Q sky130_fd_sc_hd__dfxtp_2
X_15862_ _15862_/A vssd1 vssd1 vccd1 vccd1 _18936_/D sky130_fd_sc_hd__clkbuf_1
X_17601_ _19658_/Q _16838_/A _17601_/S vssd1 vssd1 vccd1 vccd1 _17602_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14813_ _14873_/A _14813_/B _14813_/C _14813_/D vssd1 vssd1 vccd1 vccd1 _14813_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_18_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18581_ _18585_/CLK _18581_/D vssd1 vssd1 vccd1 vccd1 _18581_/Q sky130_fd_sc_hd__dfxtp_1
X_15793_ _15793_/A vssd1 vssd1 vccd1 vccd1 _15802_/S sky130_fd_sc_hd__buf_4
XFILLER_18_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16088__S _16097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17532_ _17532_/A vssd1 vssd1 vccd1 vccd1 _19627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14744_ _14875_/A vssd1 vssd1 vccd1 vccd1 _14744_/X sky130_fd_sc_hd__buf_2
X_11956_ _11956_/A _11956_/B vssd1 vssd1 vccd1 vccd1 _11956_/X sky130_fd_sc_hd__xor2_4
XFILLER_45_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13207__B1 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17463_ _17463_/A _17535_/B vssd1 vssd1 vccd1 vccd1 _17520_/A sky130_fd_sc_hd__nor2_4
X_10907_ _18851_/Q _19309_/Q _10983_/S vssd1 vssd1 vccd1 vccd1 _10907_/X sky130_fd_sc_hd__mux2_1
X_11887_ _13215_/A _11758_/X _11888_/D _18358_/Q vssd1 vssd1 vccd1 vccd1 _11887_/X
+ sky130_fd_sc_hd__a31o_1
X_14675_ _18207_/A _15959_/B vssd1 vssd1 vccd1 vccd1 _18578_/D sky130_fd_sc_hd__nor2_1
XFILLER_60_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19202_ _19427_/CLK _19202_/D vssd1 vssd1 vccd1 vccd1 _19202_/Q sky130_fd_sc_hd__dfxtp_1
X_16414_ _16414_/A vssd1 vssd1 vccd1 vccd1 _19171_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13626_ _13621_/X _13624_/X _13768_/S vssd1 vssd1 vccd1 vccd1 _13626_/X sky130_fd_sc_hd__mux2_1
X_10838_ _18591_/Q _19280_/Q _10886_/S vssd1 vssd1 vccd1 vccd1 _10838_/X sky130_fd_sc_hd__mux2_1
X_17394_ _16743_/X _19565_/Q _17402_/S vssd1 vssd1 vccd1 vccd1 _17395_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09426__A2 _09624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19133_ _19647_/CLK _19133_/D vssd1 vssd1 vccd1 vccd1 _19133_/Q sky130_fd_sc_hd__dfxtp_1
X_16345_ _16119_/X _19141_/Q _16351_/S vssd1 vssd1 vccd1 vccd1 _16346_/A sky130_fd_sc_hd__mux2_1
X_10769_ _10650_/S _10736_/Y _10768_/Y _09353_/A vssd1 vssd1 vccd1 vccd1 _10769_/Y
+ sky130_fd_sc_hd__a211oi_2
X_13557_ _13560_/A _13557_/B vssd1 vssd1 vccd1 vccd1 _13558_/A sky130_fd_sc_hd__and2_1
XFILLER_34_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15021__A _16725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12508_ _13775_/S vssd1 vssd1 vccd1 vccd1 _13742_/S sky130_fd_sc_hd__clkbuf_2
X_19064_ _19647_/CLK _19064_/D vssd1 vssd1 vccd1 vccd1 _19064_/Q sky130_fd_sc_hd__dfxtp_1
X_13488_ _13499_/A vssd1 vssd1 vccd1 vccd1 _13497_/S sky130_fd_sc_hd__buf_2
X_16276_ _16276_/A vssd1 vssd1 vccd1 vccd1 _19110_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18015_ _18027_/A _18015_/B vssd1 vssd1 vccd1 vccd1 _18015_/Y sky130_fd_sc_hd__nor2_1
X_12439_ _18380_/Q _12439_/B vssd1 vssd1 vccd1 vccd1 _12455_/B sky130_fd_sc_hd__nand2_1
XFILLER_145_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15227_ _18678_/Q _15226_/X _15233_/S vssd1 vssd1 vccd1 vccd1 _15228_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15158_ _15158_/A vssd1 vssd1 vccd1 vccd1 _18656_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11092__S1 _09538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14109_ _14126_/A _12008_/A _13975_/A _14108_/Y vssd1 vssd1 vccd1 vccd1 _14109_/X
+ sky130_fd_sc_hd__a211o_1
X_15089_ _14557_/A _11696_/Y _15092_/S vssd1 vssd1 vccd1 vccd1 _15089_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18917_ _19698_/CLK _18917_/D vssd1 vssd1 vccd1 vccd1 _18917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16787__A _16787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09650_ _19656_/Q _19073_/Q _19110_/Q _18716_/Q _11153_/A _09636_/X vssd1 vssd1 vccd1
+ vccd1 _09651_/B sky130_fd_sc_hd__mux4_1
X_18848_ _19660_/CLK _18848_/D vssd1 vssd1 vccd1 vccd1 _18848_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11427__C _12516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_clock clock vssd1 vssd1 vccd1 vccd1 clkbuf_0_clock/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__15435__A1 _15165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09581_ _10175_/A _09581_/B vssd1 vssd1 vccd1 vccd1 _09581_/Y sky130_fd_sc_hd__nor2_1
X_18779_ _19590_/CLK _18779_/D vssd1 vssd1 vccd1 vccd1 _18779_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_175_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17188__A1 _13294_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16726__S _16735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15630__S _15636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12421__A1 _13702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12154__A1_N _14559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09896__A1_N _18451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_149_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10735__A1 _10548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15077__S _15077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09917_ _09912_/Y _09915_/X _09916_/X _09919_/A vssd1 vssd1 vccd1 vccd1 _09917_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_120_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11618__B _11618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13685__A0 _14168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09848_ _09992_/A vssd1 vssd1 vccd1 vccd1 _09919_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10594__S0 _09522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09779_ _09908_/A vssd1 vssd1 vccd1 vccd1 _09905_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11810_/A _11843_/A vssd1 vssd1 vccd1 vccd1 _11844_/B sky130_fd_sc_hd__xor2_4
XFILLER_37_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12790_ _12790_/A _16847_/A _12790_/C _12790_/D vssd1 vssd1 vccd1 vccd1 _12790_/X
+ sky130_fd_sc_hd__or4_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _11741_/A _14036_/S vssd1 vssd1 vccd1 vccd1 _11785_/A sky130_fd_sc_hd__xnor2_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15540__S _15552_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17321__A _17389_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11672_ _18347_/Q _18340_/Q vssd1 vssd1 vccd1 vccd1 _11672_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _14460_/A vssd1 vssd1 vccd1 vccd1 _18501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13411_ hold3/A _13411_/B vssd1 vssd1 vccd1 vccd1 _13411_/X sky130_fd_sc_hd__or2_1
XFILLER_41_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10623_ _19637_/Q _19054_/Q _19091_/Q _18697_/Q _10605_/S _10366_/A vssd1 vssd1 vccd1
+ vccd1 _10624_/B sky130_fd_sc_hd__mux4_1
X_14391_ _14391_/A vssd1 vssd1 vccd1 vccd1 _18475_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12465__A _12465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13342_ _13045_/B _13178_/A _12749_/A _18086_/B vssd1 vssd1 vccd1 vccd1 _13342_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16130_ _16130_/A vssd1 vssd1 vccd1 vccd1 _19043_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17887__C1 _14585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10554_ _12476_/B _10554_/B vssd1 vssd1 vccd1 vccd1 _11081_/A sky130_fd_sc_hd__and2b_1
XFILLER_127_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13273_ _13273_/A _13273_/B vssd1 vssd1 vccd1 vccd1 _14859_/B sky130_fd_sc_hd__or2_1
XFILLER_6_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16061_ _16771_/A vssd1 vssd1 vccd1 vccd1 _16061_/X sky130_fd_sc_hd__clkbuf_1
X_10485_ _10239_/A _10485_/B vssd1 vssd1 vccd1 vccd1 _10485_/X sky130_fd_sc_hd__and2b_1
XFILLER_154_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12224_ _12196_/X _12220_/X _12223_/X vssd1 vssd1 vccd1 vccd1 _12224_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09774__A _10093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15012_ _15012_/A vssd1 vssd1 vccd1 vccd1 _18611_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13912__A1 _18429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10187__C1 _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19820_ _19822_/CLK _19820_/D vssd1 vssd1 vccd1 vccd1 _19820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12155_ _12155_/A _12155_/B vssd1 vssd1 vccd1 vccd1 _14192_/A sky130_fd_sc_hd__nand2_2
Xclkbuf_3_2_0_clock clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__10713__A _10713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11106_ _19416_/Q _19192_/Q _19709_/Q _19160_/Q _10230_/X _10245_/X vssd1 vssd1 vccd1
+ vccd1 _11107_/B sky130_fd_sc_hd__mux4_1
X_19751_ _19759_/CLK _19751_/D vssd1 vssd1 vccd1 vccd1 _19751_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_123_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12086_ _12086_/A _12086_/B vssd1 vssd1 vccd1 vccd1 _12089_/A sky130_fd_sc_hd__nor2_2
X_16963_ _16963_/A vssd1 vssd1 vccd1 vccd1 _19389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15715__S _15719_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18702_ _19546_/CLK _18702_/D vssd1 vssd1 vccd1 vccd1 _18702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15914_ _15914_/A vssd1 vssd1 vccd1 vccd1 _18959_/D sky130_fd_sc_hd__clkbuf_1
X_11037_ _11041_/A _11037_/B vssd1 vssd1 vccd1 vccd1 _11037_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19682_ _19682_/CLK _19682_/D vssd1 vssd1 vccd1 vccd1 _19682_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_65_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16894_ _19359_/Q _16705_/X _16902_/S vssd1 vssd1 vccd1 vccd1 _16895_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10585__S0 _10511_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18633_ _19062_/CLK _18633_/D vssd1 vssd1 vccd1 vccd1 _18633_/Q sky130_fd_sc_hd__dfxtp_2
X_15845_ _15845_/A vssd1 vssd1 vccd1 vccd1 _18928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18564_ _18564_/CLK _18564_/D vssd1 vssd1 vccd1 vccd1 _18564_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15776_ _14918_/X _18898_/Q _15780_/S vssd1 vssd1 vccd1 vccd1 _15777_/A sky130_fd_sc_hd__mux2_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12100__B1 _17241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12988_ _18310_/Q vssd1 vssd1 vccd1 vccd1 _12993_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17515_ _17515_/A vssd1 vssd1 vccd1 vccd1 _19619_/D sky130_fd_sc_hd__clkbuf_1
X_14727_ input12/X _14703_/X _14726_/X _14711_/X vssd1 vssd1 vccd1 vccd1 _16645_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10111__C1 _09988_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11939_ _11939_/A _11939_/B _14059_/B _11913_/Y vssd1 vssd1 vccd1 vccd1 _12030_/A
+ sky130_fd_sc_hd__or4b_2
X_18495_ _19693_/CLK _18495_/D vssd1 vssd1 vccd1 vccd1 _18495_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14855__A _16680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_131_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19080_/CLK sky130_fd_sc_hd__clkbuf_16
X_17446_ _16822_/X _19589_/Q _17446_/S vssd1 vssd1 vccd1 vccd1 _17447_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14658_ _14677_/A _17779_/B vssd1 vssd1 vccd1 vccd1 _14659_/A sky130_fd_sc_hd__and2_1
XANTENNA__17590__A1 _16822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13600__A0 _12011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13609_ _14126_/B _14168_/B _13681_/S vssd1 vssd1 vccd1 vccd1 _13609_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11206__A2 _11204_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17377_ _16825_/X _19558_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _17378_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14589_ _14589_/A _14589_/B vssd1 vssd1 vccd1 vccd1 _14589_/X sky130_fd_sc_hd__or2_1
X_19116_ _19630_/CLK _19116_/D vssd1 vssd1 vccd1 vccd1 _19116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16328_ _16328_/A vssd1 vssd1 vccd1 vccd1 _19133_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12094__B _19735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_146_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19597_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17377__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19047_ _19630_/CLK _19047_/D vssd1 vssd1 vccd1 vccd1 _19047_/Q sky130_fd_sc_hd__dfxtp_1
X_16259_ _16270_/A vssd1 vssd1 vccd1 vccd1 _16268_/S sky130_fd_sc_hd__buf_4
XANTENNA__16281__S _16283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11914__B1 _11970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09702_ _09172_/A _09701_/X _09184_/A vssd1 vssd1 vccd1 vccd1 _09702_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15625__S _15625_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09633_ _10422_/A vssd1 vssd1 vccd1 vccd1 _09634_/A sky130_fd_sc_hd__buf_2
XFILLER_167_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11454__A _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09564_ _09214_/A _09537_/X _09548_/X _09563_/X _09133_/A vssd1 vssd1 vccd1 vccd1
+ _09564_/X sky130_fd_sc_hd__a311o_4
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09495_ _11051_/S vssd1 vssd1 vccd1 vccd1 _10934_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16456__S _16464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15360__S _15362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14919__A0 _14918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11901__B _19737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17287__S _17291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12158__A0 _11139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10270_ _10270_/A _10270_/B vssd1 vssd1 vccd1 vccd1 _10270_/X sky130_fd_sc_hd__or2_1
XANTENNA__12732__B _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17097__A0 _16790_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__A _14431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09574__B2 _18455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13107__C1 _13102_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13960_ _13931_/A _13959_/Y _13871_/X vssd1 vssd1 vccd1 vccd1 _13960_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12911_ _12933_/C _12926_/B vssd1 vssd1 vccd1 vccd1 _12919_/C sky130_fd_sc_hd__and2_1
XFILLER_19_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13891_ _13891_/A vssd1 vssd1 vccd1 vccd1 _13970_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_46_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15630_ _18833_/Q _15542_/X _15636_/S vssd1 vssd1 vccd1 vccd1 _15631_/A sky130_fd_sc_hd__mux2_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _18263_/Q _18262_/Q _18261_/Q _12842_/D vssd1 vssd1 vccd1 vccd1 _12854_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12179__B _12180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10319__S0 _09692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _16816_/A vssd1 vssd1 vccd1 vccd1 _15561_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _18407_/Q _12768_/X _12770_/X _12772_/X vssd1 vssd1 vccd1 vccd1 _12777_/A
+ sky130_fd_sc_hd__a211o_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14675__A _18207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17300_ _19524_/Q _16715_/X _17302_/S vssd1 vssd1 vccd1 vccd1 _17301_/A sky130_fd_sc_hd__mux2_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15270__S _15278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14512_ _18524_/Q _12692_/X _14511_/X _13401_/X vssd1 vssd1 vccd1 vccd1 _18524_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18280_ _18298_/CLK _18280_/D vssd1 vssd1 vccd1 vccd1 _18280_/Q sky130_fd_sc_hd__dfxtp_1
X_11724_ _11820_/B _11721_/X _11723_/X _11676_/A vssd1 vssd1 vccd1 vccd1 _11759_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _18785_/Q _15487_/X _15504_/S vssd1 vssd1 vccd1 vccd1 _15493_/A sky130_fd_sc_hd__mux2_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17231_/A vssd1 vssd1 vccd1 vccd1 _19495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17986__A _18085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11655_ _11655_/A _11655_/B vssd1 vssd1 vccd1 vccd1 _11667_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__11811__B _13630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14443_ _18494_/Q _19732_/Q _14443_/S vssd1 vssd1 vccd1 vccd1 _14444_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_63_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19851_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12195__A _12715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10708__A _18977_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17162_ _19475_/Q _17161_/X _17172_/S vssd1 vssd1 vccd1 vccd1 _17163_/A sky130_fd_sc_hd__mux2_1
X_10606_ _09169_/A _10605_/X _09179_/A vssd1 vssd1 vccd1 vccd1 _10606_/X sky130_fd_sc_hd__a21o_1
XFILLER_167_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11586_ _13584_/C _11644_/A _13584_/D _11644_/B vssd1 vssd1 vccd1 vccd1 _11587_/C
+ sky130_fd_sc_hd__or4_1
X_14374_ _14374_/A vssd1 vssd1 vccd1 vccd1 _18469_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09801__A2 _09786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16113_ _16112_/X _19038_/Q _16113_/S vssd1 vssd1 vccd1 vccd1 _16114_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_123_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13325_ _13390_/A _18640_/Q vssd1 vssd1 vccd1 vccd1 _13325_/Y sky130_fd_sc_hd__nand2_1
X_10537_ _10530_/X _10532_/X _10534_/X _10536_/X _09245_/A vssd1 vssd1 vccd1 vccd1
+ _10537_/X sky130_fd_sc_hd__a221o_2
XFILLER_143_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17093_ _16784_/X _19447_/Q _17097_/S vssd1 vssd1 vccd1 vccd1 _17094_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16044_ _16044_/A vssd1 vssd1 vccd1 vccd1 _19016_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_78_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19727_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13256_ _13003_/B _13130_/X _12749_/A _18051_/B vssd1 vssd1 vccd1 vccd1 _13256_/X
+ sky130_fd_sc_hd__a22o_1
X_10468_ _09554_/A _10465_/X _10467_/X vssd1 vssd1 vccd1 vccd1 _10468_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12207_ _10051_/A _12328_/A _12206_/X vssd1 vssd1 vccd1 vccd1 _14216_/B sky130_fd_sc_hd__o21ai_4
XFILLER_89_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13187_ _13248_/A _18624_/Q vssd1 vssd1 vccd1 vccd1 _13187_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10399_ _19611_/Q _19449_/Q _18895_/Q _18665_/Q _10277_/S _10384_/X vssd1 vssd1 vccd1
+ vccd1 _10400_/B sky130_fd_sc_hd__mux4_1
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19803_ _19804_/CLK _19803_/D vssd1 vssd1 vccd1 vccd1 _19803_/Q sky130_fd_sc_hd__dfxtp_1
X_12138_ _12138_/A _12138_/B vssd1 vssd1 vccd1 vccd1 _12141_/A sky130_fd_sc_hd__nor2_2
XFILLER_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17995_ _19783_/Q _17997_/C _17994_/Y vssd1 vssd1 vccd1 vccd1 _19783_/D sky130_fd_sc_hd__o21a_1
XFILLER_123_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19734_ _19738_/CLK _19734_/D vssd1 vssd1 vccd1 vccd1 _19734_/Q sky130_fd_sc_hd__dfxtp_1
X_12069_ _12092_/B _12069_/B vssd1 vssd1 vccd1 vccd1 _12069_/X sky130_fd_sc_hd__and2b_1
X_16946_ _16946_/A vssd1 vssd1 vccd1 vccd1 _19381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19665_ _19687_/CLK _19665_/D vssd1 vssd1 vccd1 vccd1 _19665_/Q sky130_fd_sc_hd__dfxtp_2
X_16877_ _16877_/A vssd1 vssd1 vccd1 vccd1 _19351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18616_ _19642_/CLK _18616_/D vssd1 vssd1 vccd1 vccd1 _18616_/Q sky130_fd_sc_hd__dfxtp_1
X_15828_ _14808_/X _18921_/Q _15830_/S vssd1 vssd1 vccd1 vccd1 _15829_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_16_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19642_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19596_ _19660_/CLK _19596_/D vssd1 vssd1 vccd1 vccd1 _19596_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_48_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18547_ _19732_/CLK _18547_/D vssd1 vssd1 vccd1 vccd1 _18547_/Q sky130_fd_sc_hd__dfxtp_1
X_15759_ _15759_/A vssd1 vssd1 vccd1 vccd1 _18890_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11424__D _12537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09280_ _09280_/A vssd1 vssd1 vccd1 vccd1 _09281_/A sky130_fd_sc_hd__buf_2
X_18478_ _18519_/CLK _18478_/D vssd1 vssd1 vccd1 vccd1 _18478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17429_ _16797_/X _19581_/Q _17435_/S vssd1 vssd1 vccd1 vccd1 _17430_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10618__A _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10402__A3 _18799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17618__A2 _17617_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10353__A _10353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10549__S0 _10353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09616_ _09616_/A vssd1 vssd1 vccd1 vccd1 _09616_/X sky130_fd_sc_hd__buf_2
XFILLER_141_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14604__A2 _13106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09547_ _09172_/A _09546_/X _09184_/A vssd1 vssd1 vccd1 vccd1 _09547_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16186__S _16194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09589__A _09735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ _18978_/Q vssd1 vssd1 vccd1 vccd1 _10725_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_70_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11440_ _18550_/Q _12688_/C vssd1 vssd1 vccd1 vccd1 _11822_/B sky130_fd_sc_hd__or2_2
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10929__A1 _10996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11371_ _11736_/A _11692_/B vssd1 vssd1 vccd1 vccd1 _11371_/Y sky130_fd_sc_hd__nor2_2
XFILLER_4_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12743__A _13154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16215__A _16283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13110_ _13110_/A _13109_/X vssd1 vssd1 vccd1 vccd1 _13110_/X sky130_fd_sc_hd__or2b_1
XFILLER_152_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10322_ _09689_/X _10313_/X _10317_/X _10321_/X _09133_/A vssd1 vssd1 vccd1 vccd1
+ _10322_/X sky130_fd_sc_hd__a311o_2
X_14090_ _14320_/A _14093_/A _14088_/X _14089_/Y vssd1 vssd1 vccd1 vccd1 _14090_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13041_ _13045_/B _13045_/C _13040_/Y vssd1 vssd1 vccd1 vccd1 _18325_/D sky130_fd_sc_hd__o21a_1
XANTENNA__09547__A1 _09172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10253_ _11137_/A _12486_/A vssd1 vssd1 vccd1 vccd1 _11234_/A sky130_fd_sc_hd__or2_1
XFILLER_105_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input46_A io_ibus_inst[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ _10184_/A vssd1 vssd1 vccd1 vccd1 _10184_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16800_ _16800_/A vssd1 vssd1 vccd1 vccd1 _16800_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13574__A _13643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17780_ _17780_/A vssd1 vssd1 vccd1 vccd1 _19694_/D sky130_fd_sc_hd__clkbuf_1
X_14992_ _18450_/Q _12778_/B _14992_/S vssd1 vssd1 vccd1 vccd1 _14992_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16731_ _16731_/A vssd1 vssd1 vccd1 vccd1 _16731_/X sky130_fd_sc_hd__clkbuf_2
X_13943_ _13943_/A _13943_/B vssd1 vssd1 vccd1 vccd1 _13943_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19450_ _19551_/CLK _19450_/D vssd1 vssd1 vccd1 vccd1 _19450_/Q sky130_fd_sc_hd__dfxtp_1
X_16662_ _19281_/Q _16661_/X _16671_/S vssd1 vssd1 vccd1 vccd1 _16663_/A sky130_fd_sc_hd__mux2_1
X_13874_ _11667_/B _13827_/X _13873_/X vssd1 vssd1 vccd1 vccd1 _13874_/Y sky130_fd_sc_hd__a21oi_1
X_18401_ _18401_/CLK _18401_/D vssd1 vssd1 vccd1 vccd1 _18401_/Q sky130_fd_sc_hd__dfxtp_1
X_15613_ _15613_/A vssd1 vssd1 vccd1 vccd1 _18825_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12825_ _12844_/A _12830_/C vssd1 vssd1 vccd1 vccd1 _12825_/Y sky130_fd_sc_hd__nor2_1
X_19381_ _19543_/CLK _19381_/D vssd1 vssd1 vccd1 vccd1 _19381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16593_ _19252_/Q vssd1 vssd1 vccd1 vccd1 _16594_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_90_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18332_ _19866_/CLK _18332_/D vssd1 vssd1 vccd1 vccd1 _18332_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15544_ _15544_/A vssd1 vssd1 vccd1 vccd1 _18801_/D sky130_fd_sc_hd__clkbuf_1
X_12756_ _18642_/Q _12756_/B vssd1 vssd1 vccd1 vccd1 _12756_/X sky130_fd_sc_hd__or2_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ _19859_/CLK _18263_/D vssd1 vssd1 vccd1 vccd1 _18263_/Q sky130_fd_sc_hd__dfxtp_1
X_11707_ _19731_/Q _11752_/C vssd1 vssd1 vccd1 vccd1 _11707_/X sky130_fd_sc_hd__xor2_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15475_ _18779_/Q _15223_/X _15481_/S vssd1 vssd1 vccd1 vccd1 _15476_/A sky130_fd_sc_hd__mux2_1
X_12687_ _12661_/X _13112_/A _12780_/S vssd1 vssd1 vccd1 vccd1 _12687_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17214_ _17214_/A vssd1 vssd1 vccd1 vccd1 _19490_/D sky130_fd_sc_hd__clkbuf_1
X_14426_ _14426_/A vssd1 vssd1 vccd1 vccd1 _15087_/S sky130_fd_sc_hd__buf_2
X_18194_ _18197_/A _18194_/B vssd1 vssd1 vccd1 vccd1 _18194_/Y sky130_fd_sc_hd__nor2_1
X_11638_ _18563_/Q _11371_/Y _11535_/A _11637_/X vssd1 vssd1 vccd1 vccd1 _11638_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_129_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11968__S _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17145_ _17145_/A vssd1 vssd1 vccd1 vccd1 _19470_/D sky130_fd_sc_hd__clkbuf_1
X_14357_ _14357_/A vssd1 vssd1 vccd1 vccd1 _18463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11569_ _11729_/A vssd1 vssd1 vccd1 vccd1 _11625_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13308_ _13438_/B vssd1 vssd1 vccd1 vccd1 _13319_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17076_ _17076_/A vssd1 vssd1 vccd1 vccd1 _19439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14288_ _14323_/A _14288_/B vssd1 vssd1 vccd1 vccd1 _14288_/Y sky130_fd_sc_hd__nor2_1
X_16027_ _15055_/X _19011_/Q _16027_/S vssd1 vssd1 vccd1 vccd1 _16028_/A sky130_fd_sc_hd__mux2_1
X_13239_ _19668_/Q _12668_/X _12768_/X _18392_/Q vssd1 vssd1 vccd1 vccd1 _13240_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17978_ _19777_/Q _17979_/C _19778_/Q vssd1 vssd1 vccd1 vccd1 _17980_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__13098__A1 _18343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19717_ _19717_/CLK _19717_/D vssd1 vssd1 vccd1 vccd1 _19717_/Q sky130_fd_sc_hd__dfxtp_1
X_16929_ _16755_/X _19374_/Q _16931_/S vssd1 vssd1 vccd1 vccd1 _16930_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11144__B_N _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09710__A1 _09689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19648_ _19648_/CLK _19648_/D vssd1 vssd1 vccd1 vccd1 _19648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10951__S0 _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09401_ _10494_/A vssd1 vssd1 vccd1 vccd1 _09402_/A sky130_fd_sc_hd__buf_2
X_19579_ _19579_/CLK _19579_/D vssd1 vssd1 vccd1 vccd1 _19579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09332_ _10064_/A vssd1 vssd1 vccd1 vccd1 _09969_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09202__A _10212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09263_ _18569_/Q vssd1 vssd1 vccd1 vccd1 _14551_/A sky130_fd_sc_hd__inv_2
XFILLER_60_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09194_ _11041_/A vssd1 vssd1 vccd1 vccd1 _10875_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11033__B1 _09223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14770__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14770__B2 _14732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13089__A1 _18335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13089__B2 _13110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16909__S _16913_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15813__S _15819_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10940_ _18978_/Q vssd1 vssd1 vccd1 vccd1 _10940_/X sky130_fd_sc_hd__buf_2
XFILLER_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10871_ _10871_/A _10871_/B vssd1 vssd1 vccd1 vccd1 _10871_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12738__A _13236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_1_0_clock clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_72_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12610_ _18338_/Q _12568_/X _12546_/A _18368_/Q vssd1 vssd1 vccd1 vccd1 _12610_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _13589_/X _12450_/Y _13590_/S vssd1 vssd1 vccd1 vccd1 _13590_/X sky130_fd_sc_hd__mux2_1
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ _12566_/A _12541_/B _12541_/C vssd1 vssd1 vccd1 vccd1 _13222_/S sky130_fd_sc_hd__nor3_4
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15260_ _18687_/Q _15259_/Y _15260_/S vssd1 vssd1 vccd1 vccd1 _15261_/A sky130_fd_sc_hd__mux2_1
X_12472_ _12472_/A vssd1 vssd1 vccd1 vccd1 _12483_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14211_ _14211_/A _14319_/B vssd1 vssd1 vccd1 vccd1 _14211_/Y sky130_fd_sc_hd__nor2_1
X_11423_ _11423_/A vssd1 vssd1 vccd1 vccd1 _12686_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12473__A _12473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15191_ _16693_/A vssd1 vssd1 vccd1 vccd1 _15191_/X sky130_fd_sc_hd__buf_2
XFILLER_138_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14142_ _14142_/A _14142_/B vssd1 vssd1 vccd1 vccd1 _14142_/X sky130_fd_sc_hd__or2_1
X_11354_ _11513_/A _11514_/A _18581_/Q vssd1 vssd1 vccd1 vccd1 _11362_/A sky130_fd_sc_hd__or3_1
XFILLER_152_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12192__B _13529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10305_ _11166_/A _10305_/B vssd1 vssd1 vccd1 vccd1 _10305_/X sky130_fd_sc_hd__or2_1
XFILLER_125_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14073_ _13810_/X _13917_/X _13819_/X vssd1 vssd1 vccd1 vccd1 _14073_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_4_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18950_ _19506_/CLK _18950_/D vssd1 vssd1 vccd1 vccd1 _18950_/Q sky130_fd_sc_hd__dfxtp_1
X_11285_ _11285_/A _11285_/B vssd1 vssd1 vccd1 vccd1 _13585_/A sky130_fd_sc_hd__and2_1
XFILLER_141_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09615__S1 _10331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17901_ _17901_/A vssd1 vssd1 vccd1 vccd1 _19751_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09782__A _09782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13024_ _18320_/Q _13024_/B _13024_/C vssd1 vssd1 vccd1 vccd1 _13025_/C sky130_fd_sc_hd__and3_1
X_10236_ _10447_/A _10236_/B vssd1 vssd1 vccd1 vccd1 _10236_/Y sky130_fd_sc_hd__nor2_1
X_18881_ _19436_/CLK _18881_/D vssd1 vssd1 vccd1 vccd1 _18881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17832_ _15207_/X _19717_/Q _17838_/S vssd1 vssd1 vccd1 vccd1 _17833_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10167_ _10167_/A _10167_/B vssd1 vssd1 vccd1 vccd1 _10167_/X sky130_fd_sc_hd__or2_1
XFILLER_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17763_ _19688_/Q _17762_/X _17772_/S vssd1 vssd1 vccd1 vccd1 _17764_/A sky130_fd_sc_hd__mux2_1
X_14975_ _16816_/A vssd1 vssd1 vccd1 vccd1 _14975_/X sky130_fd_sc_hd__clkbuf_2
X_10098_ _09278_/A _10084_/X _10097_/X _09285_/A _18446_/Q vssd1 vssd1 vccd1 vccd1
+ _10098_/X sky130_fd_sc_hd__a32o_4
XANTENNA__17215__A0 _18448_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11028__S _11028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16714_ _16714_/A vssd1 vssd1 vccd1 vccd1 _19297_/D sky130_fd_sc_hd__clkbuf_1
X_19502_ _19697_/CLK _19502_/D vssd1 vssd1 vccd1 vccd1 _19502_/Q sky130_fd_sc_hd__dfxtp_1
X_13926_ _14078_/A _13924_/Y _13925_/Y _13711_/B vssd1 vssd1 vccd1 vccd1 _13926_/X
+ sky130_fd_sc_hd__a211o_1
X_17694_ _12559_/X _17692_/Y _17734_/S vssd1 vssd1 vccd1 vccd1 _17694_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19433_ _19726_/CLK _19433_/D vssd1 vssd1 vccd1 vccd1 _19433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16645_ _16645_/A vssd1 vssd1 vccd1 vccd1 _16645_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13857_ _14250_/A vssd1 vssd1 vccd1 vccd1 _14320_/A sky130_fd_sc_hd__clkbuf_2
X_12808_ _18253_/Q _12808_/B _18250_/B vssd1 vssd1 vccd1 vccd1 _12809_/C sky130_fd_sc_hd__and3_1
X_19364_ _19556_/CLK _19364_/D vssd1 vssd1 vccd1 vccd1 _19364_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13252__A1 _19669_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16576_ _16576_/A vssd1 vssd1 vccd1 vccd1 _19243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13788_ _13788_/A vssd1 vssd1 vccd1 vccd1 _13821_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18315_ _19806_/CLK _18315_/D vssd1 vssd1 vccd1 vccd1 _18315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15527_ _18796_/Q _15526_/X _15536_/S vssd1 vssd1 vccd1 vccd1 _15528_/A sky130_fd_sc_hd__mux2_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ _18290_/Q _13270_/B vssd1 vssd1 vccd1 vccd1 _12739_/X sky130_fd_sc_hd__and2_1
X_19295_ _19295_/CLK _19295_/D vssd1 vssd1 vccd1 vccd1 _19295_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18980__D _18980_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15959__A _17774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16554__S _16558_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09471__A3 _09470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18246_ _18247_/B _18247_/C _18245_/Y vssd1 vssd1 vccd1 vccd1 _19870_/D sky130_fd_sc_hd__o21a_1
X_15458_ _15458_/A vssd1 vssd1 vccd1 vccd1 _18771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14409_ _18482_/Q vssd1 vssd1 vccd1 vccd1 _14990_/A sky130_fd_sc_hd__clkbuf_2
X_18177_ _19846_/Q _18177_/B vssd1 vssd1 vccd1 vccd1 _18183_/C sky130_fd_sc_hd__and2_1
XFILLER_156_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15389_ _18742_/Q _15207_/X _15395_/S vssd1 vssd1 vccd1 vccd1 _15390_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17128_ _16835_/X _19463_/Q _17130_/S vssd1 vssd1 vccd1 vccd1 _17129_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17385__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09950_ _09927_/X _09940_/X _09949_/X _09309_/X _18449_/Q vssd1 vssd1 vccd1 vccd1
+ _12495_/C sky130_fd_sc_hd__a32o_4
X_17059_ _17059_/A vssd1 vssd1 vccd1 vccd1 _19432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09692__A _09692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09881_ _09881_/A vssd1 vssd1 vccd1 vccd1 _09881_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_112_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09931__A1 _09810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10631__A _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16729__S _16735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17206__A0 _19488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__S0 _10185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13491__A1 _13334_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10924__S0 _10919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12558__A _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11462__A _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13243__A1 _19769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09315_ _09315_/A vssd1 vssd1 vccd1 vccd1 _09621_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16464__S _16464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18182__A1 _19847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14773__A _15077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09289__D _18574_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09867__A _09867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09246_ _09246_/A vssd1 vssd1 vccd1 vccd1 _09247_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_21_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09177_ _09177_/A vssd1 vssd1 vccd1 vccd1 _10996_/A sky130_fd_sc_hd__buf_2
XFILLER_135_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11101__S0 _09449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11070_ _11070_/A _12462_/A vssd1 vssd1 vccd1 vccd1 _11254_/A sky130_fd_sc_hd__nor2_1
XFILLER_115_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10517__C1 _09314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput79 _12066_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[15] sky130_fd_sc_hd__buf_2
X_10021_ _19522_/Q _19136_/Q _19586_/Q _18742_/Q _10075_/S _09147_/A vssd1 vssd1 vccd1
+ vccd1 _10022_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09922__A1 _09217_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15109__A _15116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14259__A0 _18450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15543__S _15552_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14760_ _16654_/A vssd1 vssd1 vccd1 vccd1 _16758_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13482__A1 _12598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11972_ _12106_/A _11972_/B vssd1 vssd1 vccd1 vccd1 _11973_/B sky130_fd_sc_hd__nor2_2
XFILLER_56_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13711_ _13711_/A _13711_/B vssd1 vssd1 vccd1 vccd1 _13711_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10923_ _10923_/A vssd1 vssd1 vccd1 vccd1 _10973_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14691_ _14694_/A _14691_/B vssd1 vssd1 vccd1 vccd1 _14692_/A sky130_fd_sc_hd__and2_1
XFILLER_45_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12468__A _12468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16430_ _16430_/A _16919_/B _16919_/C vssd1 vssd1 vccd1 vccd1 _17783_/B sky130_fd_sc_hd__and3_2
XFILLER_112_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13642_ _13671_/A _12424_/A _13659_/S vssd1 vssd1 vccd1 vccd1 _13642_/X sky130_fd_sc_hd__mux2_1
X_10854_ _10850_/A _10851_/X _10853_/X _10793_/X vssd1 vssd1 vccd1 vccd1 _10854_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12037__A2 _12011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _19147_/Q _15487_/X _16369_/S vssd1 vssd1 vccd1 vccd1 _16362_/A sky130_fd_sc_hd__mux2_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13573_ _13573_/A _13573_/B _13573_/C _13573_/D vssd1 vssd1 vccd1 vccd1 _13643_/A
+ sky130_fd_sc_hd__and4_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _10785_/A vssd1 vssd1 vccd1 vccd1 _10785_/X sky130_fd_sc_hd__clkbuf_4
X_18100_ _18102_/B _18102_/C _18082_/X vssd1 vssd1 vccd1 vccd1 _18100_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10143__S1 _09867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _15312_/A vssd1 vssd1 vccd1 vccd1 _18708_/D sky130_fd_sc_hd__clkbuf_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12524_ _12603_/A vssd1 vssd1 vccd1 vccd1 _12651_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19080_ _19080_/CLK _19080_/D vssd1 vssd1 vccd1 vccd1 _19080_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16292_ _16042_/X _19117_/Q _16296_/S vssd1 vssd1 vccd1 vccd1 _16293_/A sky130_fd_sc_hd__mux2_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18031_ _19797_/Q _18031_/B _18031_/C vssd1 vssd1 vccd1 vccd1 _18033_/B sky130_fd_sc_hd__and3_1
X_15243_ _16212_/D _15242_/X _12658_/A vssd1 vssd1 vccd1 vccd1 _15243_/Y sky130_fd_sc_hd__a21oi_4
X_12455_ _18381_/Q _12455_/B vssd1 vssd1 vccd1 vccd1 _12455_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_138_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11406_ _13130_/A _12639_/A _12526_/A _11406_/D vssd1 vssd1 vccd1 vccd1 _11427_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_172_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15174_ _15174_/A vssd1 vssd1 vccd1 vccd1 _18661_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12386_ _19756_/Q _12386_/B vssd1 vssd1 vccd1 vccd1 _12388_/A sky130_fd_sc_hd__nor2_1
XFILLER_99_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14125_ _14059_/A _14124_/A _14040_/X vssd1 vssd1 vccd1 vccd1 _14125_/X sky130_fd_sc_hd__o21a_1
X_11337_ _11337_/A _11339_/B _11338_/A vssd1 vssd1 vccd1 vccd1 _11528_/B sky130_fd_sc_hd__or3_2
XFILLER_140_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18933_ _19326_/CLK _18933_/D vssd1 vssd1 vccd1 vccd1 _18933_/Q sky130_fd_sc_hd__dfxtp_1
X_14056_ _13947_/X _14055_/X _14122_/S vssd1 vssd1 vccd1 vccd1 _14056_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output77_A _12013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11268_ _11269_/B _11142_/A _10100_/A _11227_/Y vssd1 vssd1 vccd1 vccd1 _11274_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_122_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13007_ _13017_/D vssd1 vssd1 vccd1 vccd1 _13015_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10219_ _10219_/A vssd1 vssd1 vccd1 vccd1 _10219_/X sky130_fd_sc_hd__buf_2
XANTENNA__10451__A _10451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11199_ _11199_/A _12502_/A vssd1 vssd1 vccd1 vccd1 _11199_/Y sky130_fd_sc_hd__nor2_1
X_18864_ _19581_/CLK _18864_/D vssd1 vssd1 vccd1 vccd1 _18864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15961__B _17064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17815_ _17815_/A vssd1 vssd1 vccd1 vccd1 _19709_/D sky130_fd_sc_hd__clkbuf_1
X_18795_ _19543_/CLK _18795_/D vssd1 vssd1 vccd1 vccd1 _18795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15453__S _15459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17746_ _19684_/Q _17708_/X _17744_/Y _17745_/X vssd1 vssd1 vccd1 vccd1 _19684_/D
+ sky130_fd_sc_hd__o22a_1
X_14958_ _14958_/A _14958_/B _14958_/C _14958_/D vssd1 vssd1 vccd1 vccd1 _14958_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13473__A1 _13279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13909_ _14097_/A vssd1 vssd1 vccd1 vccd1 _13909_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17677_ _19672_/Q _17676_/X _17681_/S vssd1 vssd1 vccd1 vccd1 _17678_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14889_ _16793_/A vssd1 vssd1 vccd1 vccd1 _14889_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16628_ _16628_/A vssd1 vssd1 vccd1 vccd1 _19269_/D sky130_fd_sc_hd__clkbuf_1
X_19416_ _19709_/CLK _19416_/D vssd1 vssd1 vccd1 vccd1 _19416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16559_ _16559_/A vssd1 vssd1 vccd1 vccd1 _19235_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19347_ _19638_/CLK _19347_/D vssd1 vssd1 vccd1 vccd1 _19347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10134__S1 _09595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09100_ _11321_/C vssd1 vssd1 vccd1 vccd1 _11468_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09687__A _09688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19278_ _19599_/CLK _19278_/D vssd1 vssd1 vccd1 vccd1 _19278_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17911__A1 _19758_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18229_ _19864_/Q _18231_/C _12948_/X vssd1 vssd1 vccd1 vccd1 _18230_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__14725__A1 _13148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_171_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15628__S _15636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13937__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09933_ _09929_/Y _09931_/X _09932_/X _09947_/A _09892_/X vssd1 vssd1 vccd1 vccd1
+ _09940_/B sky130_fd_sc_hd__o221a_1
XANTENNA__15150__A1 _15149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17843__S _17849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09864_ _09278_/X _09854_/X _09863_/X _09285_/X _18451_/Q vssd1 vssd1 vccd1 vccd1
+ _09898_/A sky130_fd_sc_hd__a32o_4
XFILLER_112_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11172__C1 _09708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _09795_/A vssd1 vssd1 vccd1 vccd1 _10153_/S sky130_fd_sc_hd__clkbuf_4
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13464__A1 _13245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09668__B1 _09412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_96_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13216__A1 _13110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16194__S _16194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18155__A1 _19838_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10570_ _10574_/A _10570_/B vssd1 vssd1 vccd1 vccd1 _10570_/X sky130_fd_sc_hd__or2_1
XANTENNA__09597__A _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09229_ _09988_/A vssd1 vssd1 vccd1 vccd1 _09230_/A sky130_fd_sc_hd__buf_2
XFILLER_154_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09818__S1 _09875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12240_ _12240_/A _12240_/B vssd1 vssd1 vccd1 vccd1 _12241_/B sky130_fd_sc_hd__or2_1
XFILLER_135_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10202__A1 _09173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12171_ _19747_/Q _12116_/X _12167_/X _12170_/Y vssd1 vssd1 vccd1 vccd1 _17893_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17319__A _17783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12751__A _14562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11950__A1 _11082_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15141__A1 _15133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11122_ _18830_/Q _19384_/Q _19546_/Q _18798_/Q _09583_/A _10451_/A vssd1 vssd1 vccd1
+ vccd1 _11123_/B sky130_fd_sc_hd__mux4_1
XFILLER_122_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15930_ _15930_/A vssd1 vssd1 vccd1 vccd1 _18966_/D sky130_fd_sc_hd__clkbuf_1
X_11053_ _10713_/X _11050_/X _11052_/X _10797_/A vssd1 vssd1 vccd1 vccd1 _11053_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_107_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11163__C1 _09708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10004_ _10003_/B _12493_/C vssd1 vssd1 vccd1 vccd1 _10005_/B sky130_fd_sc_hd__and2b_1
X_15861_ _14986_/X _18936_/Q _15863_/S vssd1 vssd1 vccd1 vccd1 _15862_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16369__S _16369_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17600_ _17600_/A vssd1 vssd1 vccd1 vccd1 _19657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13582__A _13720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14812_ _14922_/S vssd1 vssd1 vccd1 vccd1 _14839_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_18580_ _18585_/CLK _18580_/D vssd1 vssd1 vccd1 vccd1 _18580_/Q sky130_fd_sc_hd__dfxtp_1
X_15792_ _15792_/A vssd1 vssd1 vccd1 vccd1 _18905_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17531_ _19627_/Q _16737_/X _17533_/S vssd1 vssd1 vccd1 vccd1 _17532_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17989__A _18033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14743_ _14743_/A _18461_/Q vssd1 vssd1 vccd1 vccd1 _14765_/C sky130_fd_sc_hd__and2_2
X_11955_ _11925_/A _11925_/B _11919_/A vssd1 vssd1 vccd1 vccd1 _11956_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__16893__A _16904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17462_ _17462_/A vssd1 vssd1 vccd1 vccd1 _19596_/D sky130_fd_sc_hd__clkbuf_1
X_10906_ _10906_/A _10906_/B vssd1 vssd1 vccd1 vccd1 _10906_/X sky130_fd_sc_hd__and2_1
X_14674_ input50/X _14603_/X _14643_/X _14572_/A vssd1 vssd1 vccd1 vccd1 _15959_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_72_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11886_ _11563_/X _11883_/X _11884_/Y _11885_/X vssd1 vssd1 vccd1 vccd1 _11886_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19201_ _19718_/CLK _19201_/D vssd1 vssd1 vccd1 vccd1 _19201_/Q sky130_fd_sc_hd__dfxtp_1
X_16413_ _19171_/Q _15567_/X _16413_/S vssd1 vssd1 vccd1 vccd1 _16414_/A sky130_fd_sc_hd__mux2_1
X_13625_ _13625_/A vssd1 vssd1 vccd1 vccd1 _13768_/S sky130_fd_sc_hd__clkbuf_2
X_17393_ _17461_/S vssd1 vssd1 vccd1 vccd1 _17402_/S sky130_fd_sc_hd__clkbuf_4
X_10837_ _10631_/X _10835_/Y _10836_/Y _09482_/A vssd1 vssd1 vccd1 vccd1 _10837_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_32_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19132_ _19614_/CLK _19132_/D vssd1 vssd1 vccd1 vccd1 _19132_/Q sky130_fd_sc_hd__dfxtp_1
X_16344_ _16344_/A vssd1 vssd1 vccd1 vccd1 _19140_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15302__A _15324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13556_ _13570_/B _13536_/X _13537_/A _18423_/Q vssd1 vssd1 vccd1 vccd1 _13557_/B
+ sky130_fd_sc_hd__a22o_1
X_10768_ _10788_/S _18855_/Q vssd1 vssd1 vccd1 vccd1 _10768_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12507_ _13765_/S vssd1 vssd1 vccd1 vccd1 _13775_/S sky130_fd_sc_hd__clkbuf_2
X_19063_ _19614_/CLK _19063_/D vssd1 vssd1 vccd1 vccd1 _19063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16275_ _16122_/X _19110_/Q _16279_/S vssd1 vssd1 vccd1 vccd1 _16276_/A sky130_fd_sc_hd__mux2_1
X_13487_ _13487_/A vssd1 vssd1 vccd1 vccd1 _18402_/D sky130_fd_sc_hd__clkbuf_1
X_10699_ _10724_/A vssd1 vssd1 vccd1 vccd1 _10886_/S sky130_fd_sc_hd__buf_4
X_18014_ _19790_/Q _18014_/B vssd1 vssd1 vccd1 vccd1 _18015_/B sky130_fd_sc_hd__and2_1
X_15226_ _16728_/A vssd1 vssd1 vccd1 vccd1 _15226_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12438_ _18380_/Q _12439_/B vssd1 vssd1 vccd1 vccd1 _12438_/X sky130_fd_sc_hd__or2_1
XANTENNA__15380__A1 _15194_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15448__S _15448_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15157_ _18656_/Q _15155_/X _15169_/S vssd1 vssd1 vccd1 vccd1 _15158_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12369_ _12196_/X _12367_/X _12368_/Y _11801_/X vssd1 vssd1 vccd1 vccd1 _12369_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12661__A _18335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14108_ _14250_/A _14111_/A vssd1 vssd1 vccd1 vccd1 _14108_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15088_ _15088_/A vssd1 vssd1 vccd1 vccd1 _18621_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15132__B2 _11205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17409__A0 _16768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18916_ _19597_/CLK _18916_/D vssd1 vssd1 vccd1 vccd1 _18916_/Q sky130_fd_sc_hd__dfxtp_1
X_14039_ _14178_/A vssd1 vssd1 vccd1 vccd1 _14059_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18847_ _19595_/CLK _18847_/D vssd1 vssd1 vccd1 vccd1 _18847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16279__S _16279_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09580_ _19432_/Q _19208_/Q _19725_/Q _19176_/Q _09344_/A _11189_/A vssd1 vssd1 vccd1
+ vccd1 _09581_/B sky130_fd_sc_hd__mux4_1
X_18778_ _19554_/CLK _18778_/D vssd1 vssd1 vccd1 vccd1 _18778_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_118_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17729_ _17737_/C _17728_/Y _17711_/X vssd1 vssd1 vccd1 vccd1 _17729_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_35_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15911__S _15913_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11740__A _11740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12421__A2 _14310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12555__B _12555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17838__S _17838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15371__A1 _15181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15358__S _15362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13667__A _13667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10291__S0 _09342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17573__S _17579_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09916_ _19266_/Q _19037_/Q _18968_/Q _19362_/Q _09782_/X _09783_/X vssd1 vssd1 vccd1
+ vccd1 _09916_/X sky130_fd_sc_hd__mux4_2
XANTENNA__15882__A _15950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11618__C _11688_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13685__A1 _14126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09847_ _19268_/Q _19039_/Q _18970_/Q _19364_/Q _09914_/A _09770_/X vssd1 vssd1 vccd1
+ vccd1 _09847_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09778_ _09861_/A _09778_/B vssd1 vssd1 vccd1 vccd1 _09778_/X sky130_fd_sc_hd__or2_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11448__B1 _18335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16917__S _16917_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11740_/A vssd1 vssd1 vccd1 vccd1 _14036_/S sky130_fd_sc_hd__buf_2
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10671__A1 _10605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14937__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11671_ _18352_/Q vssd1 vssd1 vccd1 vccd1 _13166_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13410_ _19789_/Q _13123_/X _13407_/X _13409_/X vssd1 vssd1 vccd1 vccd1 _13411_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_23_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10622_ _10622_/A _10622_/B vssd1 vssd1 vccd1 vccd1 _10622_/X sky130_fd_sc_hd__or2_1
XFILLER_53_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14390_ _17701_/A _18507_/Q _14395_/S vssd1 vssd1 vccd1 vccd1 _14391_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13341_ _19814_/Q vssd1 vssd1 vccd1 vccd1 _18086_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__17748__S _17762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10553_ _09274_/A _10537_/X _10552_/X _09281_/A _18436_/Q vssd1 vssd1 vccd1 vccd1
+ _10554_/B sky130_fd_sc_hd__a32o_4
XFILLER_6_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16060_ _16060_/A vssd1 vssd1 vccd1 vccd1 _19021_/D sky130_fd_sc_hd__clkbuf_1
X_13272_ _19672_/Q _13251_/X _12743_/X _18396_/Q vssd1 vssd1 vccd1 vccd1 _13273_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15362__A1 _15168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10484_ _18860_/Q _19318_/Q _10486_/S vssd1 vssd1 vccd1 vccd1 _10485_/B sky130_fd_sc_hd__mux2_1
XFILLER_6_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15011_ _15009_/X _18611_/Q _15056_/S vssd1 vssd1 vccd1 vccd1 _15012_/A sky130_fd_sc_hd__mux2_1
X_12223_ _17730_/A _12221_/Y _12272_/C _17886_/A vssd1 vssd1 vccd1 vccd1 _12223_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_108_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17049__A _17049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12481__A _12481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12154_ _14559_/A _12026_/X _12226_/A _12488_/A vssd1 vssd1 vccd1 vccd1 _12155_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10282__S0 _09342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15114__B2 _11137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17483__S _17485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11097__A _11097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ _09275_/A _11095_/X _11104_/X _09282_/A _18439_/Q vssd1 vssd1 vccd1 vccd1
+ _11130_/A sky130_fd_sc_hd__a32o_4
X_19750_ _19759_/CLK _19750_/D vssd1 vssd1 vccd1 vccd1 _19750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16962_ _16803_/X _19389_/Q _16964_/S vssd1 vssd1 vccd1 vccd1 _16963_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12085_ _12085_/A _13604_/A vssd1 vssd1 vccd1 vccd1 _12086_/B sky130_fd_sc_hd__nor2_1
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09790__A _09861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18701_ _19579_/CLK _18701_/D vssd1 vssd1 vccd1 vccd1 _18701_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11687__A0 _12462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15913_ _14879_/X _18959_/Q _15913_/S vssd1 vssd1 vccd1 vccd1 _15914_/A sky130_fd_sc_hd__mux2_1
X_11036_ _19501_/Q _19115_/Q _19565_/Q _18721_/Q _10959_/X _10960_/X vssd1 vssd1 vccd1
+ vccd1 _11037_/B sky130_fd_sc_hd__mux4_2
X_16893_ _16904_/A vssd1 vssd1 vccd1 vccd1 _16902_/S sky130_fd_sc_hd__buf_4
X_19681_ _19686_/CLK _19681_/D vssd1 vssd1 vccd1 vccd1 _19681_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_65_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18632_ _18632_/CLK _18632_/D vssd1 vssd1 vccd1 vccd1 _18632_/Q sky130_fd_sc_hd__dfxtp_2
X_15844_ _14889_/X _18928_/Q _15852_/S vssd1 vssd1 vccd1 vccd1 _15845_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18563_ _18564_/CLK _18563_/D vssd1 vssd1 vccd1 vccd1 _18563_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_18_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15775_ _15775_/A vssd1 vssd1 vccd1 vccd1 _18897_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _18309_/Q _12983_/C _12986_/Y vssd1 vssd1 vccd1 vccd1 _18309_/D sky130_fd_sc_hd__o21a_1
XANTENNA__16827__S _16839_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17514_ _19619_/Q _16712_/X _17518_/S vssd1 vssd1 vccd1 vccd1 _17515_/A sky130_fd_sc_hd__mux2_1
X_14726_ _18459_/Q _14725_/X _14923_/S vssd1 vssd1 vccd1 vccd1 _14726_/X sky130_fd_sc_hd__mux2_2
X_11938_ _11984_/A _11928_/X _11935_/X _11937_/X vssd1 vssd1 vccd1 vccd1 _17874_/B
+ sky130_fd_sc_hd__o22a_1
X_18494_ _19468_/CLK _18494_/D vssd1 vssd1 vccd1 vccd1 _18494_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17445_ _17445_/A vssd1 vssd1 vccd1 vccd1 _19588_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14657_ _14557_/A _12660_/A _14649_/X input43/X vssd1 vssd1 vccd1 vccd1 _17779_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_159_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11869_ _11870_/A _13617_/A vssd1 vssd1 vccd1 vccd1 _11871_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15050__B1 _14737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13608_ _13608_/A vssd1 vssd1 vccd1 vccd1 _14168_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__15032__A _16728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17376_ _17376_/A vssd1 vssd1 vccd1 vccd1 _17385_/S sky130_fd_sc_hd__buf_4
X_14588_ _18552_/Q _14577_/X _14587_/X _14585_/X vssd1 vssd1 vccd1 vccd1 _18552_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19115_ _19632_/CLK _19115_/D vssd1 vssd1 vccd1 vccd1 _19115_/Q sky130_fd_sc_hd__dfxtp_1
X_16327_ _16093_/X _19133_/Q _16329_/S vssd1 vssd1 vccd1 vccd1 _16328_/A sky130_fd_sc_hd__mux2_1
X_13539_ _13542_/A _13539_/B vssd1 vssd1 vccd1 vccd1 _13540_/A sky130_fd_sc_hd__and2_1
XFILLER_146_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12094__C _19743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19046_ _19632_/CLK _19046_/D vssd1 vssd1 vccd1 vccd1 _19046_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09965__A _09969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16258_ _16258_/A vssd1 vssd1 vccd1 vccd1 _19102_/D sky130_fd_sc_hd__clkbuf_1
X_15209_ _15209_/A vssd1 vssd1 vccd1 vccd1 _18672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16189_ _16189_/A vssd1 vssd1 vccd1 vccd1 _19067_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15105__A1 _18629_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15105__B2 _10554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__A2 _18427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09701_ _18875_/Q _19333_/Q _09701_/S vssd1 vssd1 vccd1 vccd1 _09701_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09966__S0 _09803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15207__A _16709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09632_ _09632_/A vssd1 vssd1 vccd1 vccd1 _11153_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__14111__A _14111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09205__A _09861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09563_ _09772_/A _09556_/X _09561_/X _09562_/X vssd1 vssd1 vccd1 vccd1 _09563_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15641__S _15647_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09494_ _18977_/Q vssd1 vssd1 vccd1 vccd1 _11051_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_51_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17568__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14781__A _16661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09875__A _09875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10169__B1 _09230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09574__A2 _09564_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09957__S0 _09866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12910_ _18282_/Q _18281_/Q _18280_/Q _12910_/D vssd1 vssd1 vccd1 vccd1 _12926_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_24_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13890_ _13886_/X _13889_/X _14085_/S vssd1 vssd1 vccd1 vccd1 _13890_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12841_ _12851_/A _12841_/B _12841_/C vssd1 vssd1 vccd1 vccd1 _18262_/D sky130_fd_sc_hd__nor3_1
XFILLER_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14083__A1 _11956_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10319__S1 _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _15560_/A vssd1 vssd1 vccd1 vccd1 _18806_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17332__A _17389_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _19683_/Q _12737_/A _13203_/A _19493_/Q vssd1 vssd1 vccd1 vccd1 _12772_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13830__A1 _11022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14675__B _15959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14511_/A _14519_/B vssd1 vssd1 vccd1 vccd1 _14511_/X sky130_fd_sc_hd__or2_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11723_/A _11723_/B _11723_/C vssd1 vssd1 vccd1 vccd1 _11723_/X sky130_fd_sc_hd__and3_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15491_ _15590_/S vssd1 vssd1 vccd1 vccd1 _15504_/S sky130_fd_sc_hd__buf_2
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17230_ _19495_/Q _17229_/X _17239_/S vssd1 vssd1 vccd1 vccd1 _17231_/A sky130_fd_sc_hd__mux2_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _14442_/A vssd1 vssd1 vccd1 vccd1 _18493_/D sky130_fd_sc_hd__clkbuf_1
X_11654_ _12511_/A _11623_/B _11621_/X vssd1 vssd1 vccd1 vccd1 _11655_/B sky130_fd_sc_hd__a21o_2
XFILLER_80_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17161_ _18432_/Q _13212_/X _17167_/S vssd1 vssd1 vccd1 vccd1 _17161_/X sky130_fd_sc_hd__mux2_1
X_10605_ _18857_/Q _19315_/Q _10605_/S vssd1 vssd1 vccd1 vccd1 _10605_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14373_ _17662_/A _18501_/Q _14381_/S vssd1 vssd1 vccd1 vccd1 _14374_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11585_ _11585_/A _11585_/B _11642_/C _11585_/D vssd1 vssd1 vccd1 vccd1 _11644_/B
+ sky130_fd_sc_hd__nor4_2
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16112_ _16822_/A vssd1 vssd1 vccd1 vccd1 _16112_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09801__A3 _09800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13324_ _13324_/A vssd1 vssd1 vccd1 vccd1 _13390_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17092_ _17092_/A vssd1 vssd1 vccd1 vccd1 _19446_/D sky130_fd_sc_hd__clkbuf_1
X_10536_ _09549_/A _10535_/X _09225_/A vssd1 vssd1 vccd1 vccd1 _10536_/X sky130_fd_sc_hd__o21a_1
XFILLER_155_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16043_ _16042_/X _19016_/Q _16049_/S vssd1 vssd1 vccd1 vccd1 _16044_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13255_ _19802_/Q vssd1 vssd1 vccd1 vccd1 _18051_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__10724__A _10724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10467_ _09170_/A _10466_/X _09454_/A vssd1 vssd1 vccd1 vccd1 _10467_/X sky130_fd_sc_hd__a21o_1
XFILLER_142_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12206_ _18511_/Q _12259_/B _12259_/C vssd1 vssd1 vccd1 vccd1 _12206_/X sky130_fd_sc_hd__or3_1
XFILLER_124_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13186_ _13324_/A vssd1 vssd1 vccd1 vccd1 _13248_/A sky130_fd_sc_hd__clkbuf_2
X_10398_ _09315_/A _10386_/Y _10391_/X _10394_/Y _10397_/Y vssd1 vssd1 vccd1 vccd1
+ _10398_/X sky130_fd_sc_hd__o32a_1
XFILLER_9_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19802_ _19806_/CLK _19802_/D vssd1 vssd1 vccd1 vccd1 _19802_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15726__S _15730_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12137_ _12137_/A _13596_/A vssd1 vssd1 vccd1 vccd1 _12138_/B sky130_fd_sc_hd__nor2_1
XFILLER_97_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17994_ _19783_/Q _17997_/C _17993_/X vssd1 vssd1 vccd1 vccd1 _17994_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_96_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19733_ _19733_/CLK _19733_/D vssd1 vssd1 vccd1 vccd1 _19733_/Q sky130_fd_sc_hd__dfxtp_4
X_12068_ _12043_/A _12067_/B _12067_/D _19743_/Q vssd1 vssd1 vccd1 vccd1 _12069_/B
+ sky130_fd_sc_hd__a31o_1
X_16945_ _16777_/X _19381_/Q _16953_/S vssd1 vssd1 vccd1 vccd1 _16946_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12321__A1 _17711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ _11065_/A _11019_/B vssd1 vssd1 vccd1 vccd1 _11019_/X sky130_fd_sc_hd__or2_1
X_19664_ _19687_/CLK _19664_/D vssd1 vssd1 vccd1 vccd1 _19664_/Q sky130_fd_sc_hd__dfxtp_2
X_16876_ _19351_/Q _16680_/X _16880_/S vssd1 vssd1 vccd1 vccd1 _16877_/A sky130_fd_sc_hd__mux2_1
X_18615_ _19724_/CLK _18615_/D vssd1 vssd1 vccd1 vccd1 _18615_/Q sky130_fd_sc_hd__dfxtp_1
X_15827_ _15827_/A vssd1 vssd1 vccd1 vccd1 _18920_/D sky130_fd_sc_hd__clkbuf_1
X_19595_ _19595_/CLK _19595_/D vssd1 vssd1 vccd1 vccd1 _19595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14866__A _16683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18546_ _19481_/CLK _18546_/D vssd1 vssd1 vccd1 vccd1 _18546_/Q sky130_fd_sc_hd__dfxtp_1
X_15758_ _14821_/X _18890_/Q _15758_/S vssd1 vssd1 vccd1 vccd1 _15759_/A sky130_fd_sc_hd__mux2_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14709_ _19080_/Q vssd1 vssd1 vccd1 vccd1 _14903_/A sky130_fd_sc_hd__inv_2
XANTENNA__12386__A _19756_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15689_ _18859_/Q _15522_/X _15697_/S vssd1 vssd1 vccd1 vccd1 _15690_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18477_ _18510_/CLK _18477_/D vssd1 vssd1 vccd1 vccd1 _18477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17428_ _17428_/A vssd1 vssd1 vccd1 vccd1 _19580_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16292__S _16296_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17359_ _16800_/X _19550_/Q _17363_/S vssd1 vssd1 vccd1 vccd1 _17360_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11805__A2_N _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09695__A _09695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14129__A2 _14126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19029_ _19612_/CLK _19029_/D vssd1 vssd1 vccd1 vccd1 _19029_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_146_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10634__A _10634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10246__S0 _10279_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15636__S _15636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10549__S1 _10548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17851__S _17853_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09615_ _19658_/Q _19075_/Q _19112_/Q _18718_/Q _09729_/S _10331_/A vssd1 vssd1 vccd1
+ vccd1 _09615_/X sky130_fd_sc_hd__mux4_2
XFILLER_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15371__S _15373_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ _18878_/Q _19336_/Q _09793_/A vssd1 vssd1 vccd1 vccd1 _09546_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_0_0_clock_A clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ _09522_/A vssd1 vssd1 vccd1 vccd1 _10389_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_54_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_192_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19223_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17298__S _17302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11370_ _11736_/B vssd1 vssd1 vccd1 vccd1 _11692_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10321_ _11166_/A _10318_/X _10320_/X _09562_/X vssd1 vssd1 vccd1 vccd1 _10321_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13040_ _13045_/B _13045_/C _13011_/X vssd1 vssd1 vccd1 vccd1 _13040_/Y sky130_fd_sc_hd__a21oi_1
X_10252_ _18443_/Q _09308_/A _09429_/A _10251_/X vssd1 vssd1 vccd1 vccd1 _12486_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15546__S _15552_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10183_ _18867_/Q _19325_/Q _11188_/S vssd1 vssd1 vccd1 vccd1 _10184_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_130_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19081_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_132_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input39_A io_ibus_inst[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14991_ _14990_/A _15002_/C _14815_/A vssd1 vssd1 vccd1 vccd1 _14991_/X sky130_fd_sc_hd__o21a_1
XFILLER_94_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13942_ _13942_/A vssd1 vssd1 vccd1 vccd1 _13943_/A sky130_fd_sc_hd__clkbuf_2
X_16730_ _16730_/A vssd1 vssd1 vccd1 vccd1 _19302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_145_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19697_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_46_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16661_ _16661_/A vssd1 vssd1 vccd1 vccd1 _16661_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13873_ _14173_/A vssd1 vssd1 vccd1 vccd1 _13873_/X sky130_fd_sc_hd__buf_4
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18400_ _18401_/CLK _18400_/D vssd1 vssd1 vccd1 vccd1 _18400_/Q sky130_fd_sc_hd__dfxtp_1
X_15612_ _18825_/Q _15516_/X _15614_/S vssd1 vssd1 vccd1 vccd1 _15613_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12824_ _12832_/D vssd1 vssd1 vccd1 vccd1 _12830_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19380_ _19541_/CLK _19380_/D vssd1 vssd1 vccd1 vccd1 _19380_/Q sky130_fd_sc_hd__dfxtp_1
X_16592_ _16592_/A vssd1 vssd1 vccd1 vccd1 _19251_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18331_ _19866_/CLK _18331_/D vssd1 vssd1 vccd1 vccd1 _18331_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11822__B _11822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15543_ _18801_/Q _15542_/X _15552_/S vssd1 vssd1 vccd1 vccd1 _15544_/A sky130_fd_sc_hd__mux2_1
X_12755_ _19847_/Q _12736_/X _12745_/X _12750_/X _12754_/X vssd1 vssd1 vccd1 vccd1
+ _12756_/B sky130_fd_sc_hd__a2111o_2
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15005__A0 _18451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10719__A _10724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18262_ _19855_/CLK _18262_/D vssd1 vssd1 vccd1 vccd1 _18262_/Q sky130_fd_sc_hd__dfxtp_1
X_11706_ _14431_/B vssd1 vssd1 vccd1 vccd1 _11706_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _15474_/A vssd1 vssd1 vccd1 vccd1 _18778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16753__A0 _16752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12686_ _12686_/A _12791_/A _12791_/B _13108_/B vssd1 vssd1 vccd1 vccd1 _12780_/S
+ sky130_fd_sc_hd__nor4_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17213_ _19490_/Q _17212_/X _17223_/S vssd1 vssd1 vccd1 vccd1 _17214_/A sky130_fd_sc_hd__mux2_1
X_14425_ _14425_/A vssd1 vssd1 vccd1 vccd1 _18487_/D sky130_fd_sc_hd__clkbuf_1
X_18193_ _19852_/Q _18196_/C vssd1 vssd1 vccd1 vccd1 _18194_/B sky130_fd_sc_hd__and2_1
X_11637_ _11736_/A _11692_/B _11637_/C vssd1 vssd1 vccd1 vccd1 _11637_/X sky130_fd_sc_hd__or3_1
XANTENNA__17001__S _17003_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17144_ _19470_/Q _17143_/X _17155_/S vssd1 vssd1 vccd1 vccd1 _17145_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10476__S0 _09631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14356_ _17632_/A _18495_/Q _14367_/S vssd1 vssd1 vccd1 vccd1 _14357_/A sky130_fd_sc_hd__mux2_1
X_11568_ input66/X _12715_/A vssd1 vssd1 vccd1 vccd1 _11729_/A sky130_fd_sc_hd__nand2_1
XFILLER_156_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13307_ _13297_/X _13298_/Y _13305_/X _13306_/X _18634_/Q vssd1 vssd1 vccd1 vccd1
+ _13307_/X sky130_fd_sc_hd__a32o_4
XANTENNA__10250__C1 _09393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17075_ _16758_/X _19439_/Q _17075_/S vssd1 vssd1 vccd1 vccd1 _17076_/A sky130_fd_sc_hd__mux2_1
X_10519_ _19511_/Q _19125_/Q _19575_/Q _18731_/Q _10500_/X _10238_/A vssd1 vssd1 vccd1
+ vccd1 _10520_/B sky130_fd_sc_hd__mux4_2
XFILLER_6_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14287_ _14289_/A _14289_/B vssd1 vssd1 vccd1 vccd1 _14288_/B sky130_fd_sc_hd__and2_1
X_11499_ _11551_/A _11528_/A _11664_/D vssd1 vssd1 vccd1 vccd1 _11511_/C sky130_fd_sc_hd__or3_1
XFILLER_115_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16026_ _16026_/A vssd1 vssd1 vccd1 vccd1 _19010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13238_ _19478_/Q _13235_/X _13236_/X _13246_/A _13237_/X vssd1 vssd1 vccd1 vccd1
+ _13240_/A sky130_fd_sc_hd__a221o_1
XFILLER_108_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10228__S0 _09583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12542__A1 _19675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13169_ _13112_/A _13183_/B _14673_/A vssd1 vssd1 vccd1 vccd1 _13169_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16141__A _16209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17977_ _19777_/Q _17979_/C _17976_/Y vssd1 vssd1 vccd1 vccd1 _19777_/D sky130_fd_sc_hd__o21a_1
XANTENNA__13098__A2 _12731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14295__A1 _18453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14295__B2 _14294_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19716_ _19716_/CLK _19716_/D vssd1 vssd1 vccd1 vccd1 _19716_/Q sky130_fd_sc_hd__dfxtp_1
X_16928_ _16928_/A vssd1 vssd1 vccd1 vccd1 _19373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10856__B2 _18431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19647_ _19647_/CLK _19647_/D vssd1 vssd1 vccd1 vccd1 _19647_/Q sky130_fd_sc_hd__dfxtp_1
X_16859_ _16859_/A vssd1 vssd1 vccd1 vccd1 _19343_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14596__A _14612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09400_ _10589_/A vssd1 vssd1 vccd1 vccd1 _10494_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10951__S1 _10726_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19578_ _19709_/CLK _19578_/D vssd1 vssd1 vccd1 vccd1 _19578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09331_ _10140_/A vssd1 vssd1 vccd1 vccd1 _10064_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11732__B _13996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18529_ _18618_/CLK _18529_/D vssd1 vssd1 vccd1 vccd1 _18529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ _18570_/Q _16138_/A _09259_/X _09260_/Y _16212_/C vssd1 vssd1 vccd1 vccd1
+ _11368_/B sky130_fd_sc_hd__o221a_1
XFILLER_166_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09193_ _10928_/A vssd1 vssd1 vccd1 vccd1 _11041_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11033__A1 _10956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_62_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19833_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16197__S _16205_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_166_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10870_ _18822_/Q _19376_/Q _19538_/Q _18790_/Q _10664_/S _10365_/A vssd1 vssd1 vccd1
+ vccd1 _10871_/B sky130_fd_sc_hd__mux4_2
XFILLER_83_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_77_clock clkbuf_opt_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19660_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _10219_/A vssd1 vssd1 vccd1 vccd1 _09529_/X sky130_fd_sc_hd__clkbuf_4
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _12540_/A _12540_/B vssd1 vssd1 vccd1 vccd1 _12541_/C sky130_fd_sc_hd__nand2_1
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09560__S1 _09642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12471_ _13526_/A _12471_/B _12471_/C vssd1 vssd1 vccd1 vccd1 _12472_/A sky130_fd_sc_hd__or3_4
XANTENNA__16226__A _16283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14210_ _14210_/A vssd1 vssd1 vccd1 vccd1 _18446_/D sky130_fd_sc_hd__clkbuf_1
X_11422_ _12533_/A _12540_/A _12533_/B vssd1 vssd1 vccd1 vccd1 _12530_/A sky130_fd_sc_hd__or3b_1
XANTENNA__12221__B1 _18371_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15190_ _15190_/A vssd1 vssd1 vccd1 vccd1 _18666_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12772__A1 _19683_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10378__A3 _18799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14141_ _13714_/X _14142_/B _14139_/X _14140_/X vssd1 vssd1 vccd1 vccd1 _14141_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_11353_ _11598_/B _11476_/B vssd1 vssd1 vccd1 vccd1 _11360_/C sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_15_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19581_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_153_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10304_ _19644_/Q _19061_/Q _19098_/Q _18704_/Q _09553_/X _09555_/X vssd1 vssd1 vccd1
+ vccd1 _10305_/B sky130_fd_sc_hd__mux4_1
X_14072_ _13919_/X _14071_/X _14086_/S vssd1 vssd1 vccd1 vccd1 _14072_/X sky130_fd_sc_hd__mux2_1
X_11284_ _14545_/A _11284_/B _11284_/C _13568_/B vssd1 vssd1 vccd1 vccd1 _11284_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_106_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17900_ _17909_/A _17900_/B vssd1 vssd1 vccd1 vccd1 _17901_/A sky130_fd_sc_hd__and2_1
X_13023_ _13024_/B _13024_/C _18320_/Q vssd1 vssd1 vccd1 vccd1 _13025_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__15276__S _15278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10235_ _19260_/Q _19031_/Q _18962_/Q _19356_/Q _10224_/X _09486_/X vssd1 vssd1 vccd1
+ vccd1 _10236_/B sky130_fd_sc_hd__mux4_2
X_18880_ _19648_/CLK _18880_/D vssd1 vssd1 vccd1 vccd1 _18880_/Q sky130_fd_sc_hd__dfxtp_1
X_17831_ _17831_/A vssd1 vssd1 vccd1 vccd1 _19716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10166_ _19615_/Q _19453_/Q _18899_/Q _18669_/Q _10200_/S _09979_/A vssd1 vssd1 vccd1
+ vccd1 _10167_/B sky130_fd_sc_hd__mux4_1
X_17762_ _13412_/X _17761_/Y _17762_/S vssd1 vssd1 vccd1 vccd1 _17762_/X sky130_fd_sc_hd__mux2_1
X_14974_ _16712_/A vssd1 vssd1 vccd1 vccd1 _16816_/A sky130_fd_sc_hd__clkbuf_2
X_10097_ _10089_/X _10091_/X _10093_/X _10096_/X _09249_/A vssd1 vssd1 vccd1 vccd1
+ _10097_/X sky130_fd_sc_hd__a221o_1
XFILLER_59_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17215__A1 _13346_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19501_ _19697_/CLK _19501_/D vssd1 vssd1 vccd1 vccd1 _19501_/Q sky130_fd_sc_hd__dfxtp_1
X_16713_ _19297_/Q _16712_/X _16719_/S vssd1 vssd1 vccd1 vccd1 _16714_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13925_ _13999_/S _13925_/B vssd1 vssd1 vccd1 vccd1 _13925_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17693_ _17693_/A vssd1 vssd1 vccd1 vccd1 _17734_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_48_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19432_ _19725_/CLK _19432_/D vssd1 vssd1 vccd1 vccd1 _19432_/Q sky130_fd_sc_hd__dfxtp_1
X_16644_ _16644_/A vssd1 vssd1 vccd1 vccd1 _19275_/D sky130_fd_sc_hd__clkbuf_1
X_13856_ _13856_/A vssd1 vssd1 vccd1 vccd1 _13862_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12807_ _12808_/B _18250_/B _18253_/Q vssd1 vssd1 vccd1 vccd1 _12809_/B sky130_fd_sc_hd__a21oi_1
XFILLER_90_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19363_ _19589_/CLK _19363_/D vssd1 vssd1 vccd1 vccd1 _19363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16575_ _19243_/Q vssd1 vssd1 vccd1 vccd1 _16576_/A sky130_fd_sc_hd__clkbuf_1
X_13787_ _14037_/A vssd1 vssd1 vccd1 vccd1 _13788_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10999_ _10992_/Y _10994_/Y _10996_/Y _10998_/Y _19695_/Q vssd1 vssd1 vccd1 vccd1
+ _10999_/X sky130_fd_sc_hd__o221a_1
X_18314_ _19798_/CLK _18314_/D vssd1 vssd1 vccd1 vccd1 _18314_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17520__A _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12738_ _13236_/A vssd1 vssd1 vccd1 vccd1 _13115_/A sky130_fd_sc_hd__buf_2
X_15526_ _16781_/A vssd1 vssd1 vccd1 vccd1 _15526_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10697__S0 _11050_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19294_ _19648_/CLK _19294_/D vssd1 vssd1 vccd1 vccd1 _19294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15959__B _15959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18245_ _18247_/B _18247_/C _12844_/A vssd1 vssd1 vccd1 vccd1 _18245_/Y sky130_fd_sc_hd__a21oi_1
X_15457_ _18771_/Q _15197_/X _15459_/S vssd1 vssd1 vccd1 vccd1 _15458_/A sky130_fd_sc_hd__mux2_1
X_12669_ _12669_/A vssd1 vssd1 vccd1 vccd1 _13235_/A sky130_fd_sc_hd__buf_2
XFILLER_30_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14408_ _14408_/A vssd1 vssd1 vccd1 vccd1 _18481_/D sky130_fd_sc_hd__clkbuf_1
X_18176_ _18249_/A _18176_/B _18177_/B vssd1 vssd1 vccd1 vccd1 _19845_/D sky130_fd_sc_hd__nor3_1
XFILLER_129_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15388_ _15388_/A vssd1 vssd1 vccd1 vccd1 _18741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11420__D1 _12603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14339_ _18457_/Q _14120_/X _14338_/X vssd1 vssd1 vccd1 vccd1 _18457_/D sky130_fd_sc_hd__o21a_1
X_17127_ _17127_/A vssd1 vssd1 vccd1 vccd1 _19462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17058_ _19432_/Q _16734_/X _17058_/S vssd1 vssd1 vccd1 vccd1 _17059_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16009_ _16009_/A vssd1 vssd1 vccd1 vccd1 _19002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09880_ _09880_/A vssd1 vssd1 vccd1 vccd1 _09881_/A sky130_fd_sc_hd__clkbuf_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10526__B1 _09314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10621__S0 _10353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10924__S1 _10920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09213__A _09689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11462__B _13532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09314_ _09314_/A vssd1 vssd1 vccd1 vccd1 _09315_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10688__S0 _10669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09245_ _09245_/A vssd1 vssd1 vccd1 vccd1 _09246_/A sky130_fd_sc_hd__buf_4
XFILLER_166_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12574__A _17895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09176_ _10923_/A vssd1 vssd1 vccd1 vccd1 _09177_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11101__S1 _09538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16480__S _16486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10094__A _10094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_92_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10020_ _10020_/A _10020_/B vssd1 vssd1 vccd1 vccd1 _10020_/X sky130_fd_sc_hd__or2_1
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14259__A1 _14258_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10033__S _10033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11971_ _12030_/A _14075_/B vssd1 vssd1 vccd1 vccd1 _11972_/B sky130_fd_sc_hd__nor2_1
XFILLER_91_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09686__B2 _09685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13710_ _14312_/A vssd1 vssd1 vccd1 vccd1 _13806_/A sky130_fd_sc_hd__buf_2
X_10922_ _11026_/A _10922_/B vssd1 vssd1 vccd1 vccd1 _10922_/X sky130_fd_sc_hd__or2_1
XANTENNA__15125__A _15125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14690_ _14584_/A _14648_/X _14680_/X input55/X vssd1 vssd1 vccd1 vccd1 _14691_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13641_ _13635_/X _13638_/X _13743_/S vssd1 vssd1 vccd1 vccd1 _13641_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10853_ _10950_/A _10853_/B vssd1 vssd1 vccd1 vccd1 _10853_/X sky130_fd_sc_hd__or2_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16360_ _16428_/S vssd1 vssd1 vccd1 vccd1 _16369_/S sky130_fd_sc_hd__clkbuf_4
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ _13572_/A _13572_/B _13572_/C vssd1 vssd1 vccd1 vccd1 _13573_/D sky130_fd_sc_hd__and3_1
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10784_ _10691_/X _12469_/A _11252_/A vssd1 vssd1 vccd1 vccd1 _11248_/A sky130_fd_sc_hd__o21ai_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _18708_/Q _15200_/X _15311_/S vssd1 vssd1 vccd1 vccd1 _15312_/A sky130_fd_sc_hd__mux2_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _18319_/Q vssd1 vssd1 vccd1 vccd1 _13024_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ _16291_/A vssd1 vssd1 vccd1 vccd1 _19116_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12484__A _12505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15242_ _15242_/A _15242_/B _15242_/C _15242_/D vssd1 vssd1 vccd1 vccd1 _15242_/X
+ sky130_fd_sc_hd__or4_1
X_18030_ _18031_/B _18031_/C _18029_/Y vssd1 vssd1 vccd1 vccd1 _19796_/D sky130_fd_sc_hd__o21a_1
XFILLER_9_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12454_ _11980_/A _12452_/X _12453_/X _17711_/A vssd1 vssd1 vccd1 vccd1 _12454_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12745__A1 _19682_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11405_ _11423_/A _11412_/A _12747_/C vssd1 vssd1 vccd1 vccd1 _11406_/D sky130_fd_sc_hd__nor3_2
X_15173_ _18661_/Q _15171_/X _15185_/S vssd1 vssd1 vccd1 vccd1 _15174_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12385_ _12385_/A _12385_/B vssd1 vssd1 vccd1 vccd1 _12385_/X sky130_fd_sc_hd__xor2_4
XFILLER_125_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14124_ _14124_/A _14126_/B vssd1 vssd1 vccd1 vccd1 _14128_/B sky130_fd_sc_hd__and2_1
XANTENNA__09793__A _09793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11336_ _18560_/Q _18559_/Q _18558_/Q vssd1 vssd1 vccd1 vccd1 _11338_/A sky130_fd_sc_hd__or3b_1
XANTENNA__14498__A1 _19757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18932_ _19326_/CLK _18932_/D vssd1 vssd1 vccd1 vccd1 _18932_/Q sky130_fd_sc_hd__dfxtp_1
X_14055_ _13841_/X _13846_/A _14121_/S vssd1 vssd1 vccd1 vccd1 _14055_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10732__A _10732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11267_ _11227_/Y _11228_/X _11231_/X _11233_/Y _11266_/X vssd1 vssd1 vccd1 vccd1
+ _11267_/X sky130_fd_sc_hd__a2111o_1
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13006_ _18314_/Q _18313_/Q _18315_/Q _13006_/D vssd1 vssd1 vccd1 vccd1 _13017_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_79_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10218_ _09277_/A _10208_/X _10217_/X _09284_/A _18443_/Q vssd1 vssd1 vccd1 vccd1
+ _11137_/A sky130_fd_sc_hd__a32o_4
X_18863_ _19640_/CLK _18863_/D vssd1 vssd1 vccd1 vccd1 _18863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11198_ _11199_/A _12502_/A vssd1 vssd1 vccd1 vccd1 _11198_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15734__S _15734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17814_ _15181_/X _19709_/Q _17816_/S vssd1 vssd1 vccd1 vccd1 _17815_/A sky130_fd_sc_hd__mux2_1
X_10149_ _09430_/X _10138_/X _10147_/X _09625_/X _10148_/Y vssd1 vssd1 vccd1 vccd1
+ _12488_/A sky130_fd_sc_hd__o32a_4
X_18794_ _19639_/CLK _18794_/D vssd1 vssd1 vccd1 vccd1 _18794_/Q sky130_fd_sc_hd__dfxtp_1
X_17745_ _17730_/X _13364_/X _17724_/X vssd1 vssd1 vccd1 vccd1 _17745_/X sky130_fd_sc_hd__a21bo_1
XFILLER_48_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09677__A1 _10329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14957_ _14979_/C _14957_/B vssd1 vssd1 vccd1 vccd1 _14957_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12659__A _14648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13908_ _13931_/A _13908_/B _13908_/C vssd1 vssd1 vccd1 vccd1 _13908_/X sky130_fd_sc_hd__or3_1
X_17676_ _13279_/X _17675_/Y _17686_/S vssd1 vssd1 vccd1 vccd1 _17676_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14888_ _16689_/A vssd1 vssd1 vccd1 vccd1 _16793_/A sky130_fd_sc_hd__clkbuf_2
X_19415_ _19708_/CLK _19415_/D vssd1 vssd1 vccd1 vccd1 _19415_/Q sky130_fd_sc_hd__dfxtp_1
X_16627_ _19269_/Q vssd1 vssd1 vccd1 vccd1 _16628_/A sky130_fd_sc_hd__clkbuf_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13839_ _13680_/X _13690_/X _13839_/S vssd1 vssd1 vccd1 vccd1 _13839_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16565__S _16569_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19346_ _19506_/CLK _19346_/D vssd1 vssd1 vccd1 vccd1 _19346_/Q sky130_fd_sc_hd__dfxtp_1
X_16558_ _19235_/Q _15567_/X _16558_/S vssd1 vssd1 vccd1 vccd1 _16559_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15509_ _15509_/A vssd1 vssd1 vccd1 vccd1 _18790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19277_ _19599_/CLK _19277_/D vssd1 vssd1 vccd1 vccd1 _19277_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09687__B _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16175__A1 _19061_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16489_ _16115_/X _19204_/Q _16497_/S vssd1 vssd1 vccd1 vccd1 _16490_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14186__A0 _18444_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18228_ _19864_/Q _18231_/C vssd1 vssd1 vccd1 vccd1 _18230_/A sky130_fd_sc_hd__and2_1
XFILLER_30_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17396__S _17402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15909__S _15913_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18159_ _18159_/A _18164_/C vssd1 vssd1 vccd1 vccd1 _18159_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_114_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13523__C_N _14568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10842__S0 _10648_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14641__A1_N input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09932_ _19266_/Q _19037_/Q _18968_/Q _19362_/Q _09874_/S _09869_/X vssd1 vssd1 vccd1
+ vccd1 _09932_/X sky130_fd_sc_hd__mux4_2
XFILLER_131_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09863_ _09217_/X _09856_/X _09858_/X _09862_/X _09249_/X vssd1 vssd1 vccd1 vccd1
+ _09863_/X sky130_fd_sc_hd__a311o_2
XFILLER_113_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09794_/A vssd1 vssd1 vccd1 vccd1 _09795_/A sky130_fd_sc_hd__buf_4
XFILLER_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16938__A0 _16768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_39_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10435__C1 _09246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09228_ _09708_/A vssd1 vssd1 vccd1 vccd1 _09988_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12727__B2 _18631_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15819__S _15819_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09159_ _11156_/S vssd1 vssd1 vccd1 vccd1 _10154_/S sky130_fd_sc_hd__buf_2
XFILLER_147_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14723__S _14762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12170_ _12091_/A _12168_/Y _12222_/C _11859_/X vssd1 vssd1 vccd1 vccd1 _12170_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_123_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11121_ _10226_/A _11120_/X _10219_/X vssd1 vssd1 vccd1 vccd1 _11121_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_1_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11052_ _10713_/A _11052_/B vssd1 vssd1 vccd1 vccd1 _11052_/X sky130_fd_sc_hd__and2b_1
XFILLER_77_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10003_ _12493_/C _10003_/B vssd1 vssd1 vccd1 vccd1 _11272_/A sky130_fd_sc_hd__and2b_1
X_15860_ _15860_/A vssd1 vssd1 vccd1 vccd1 _18935_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input21_A io_dbus_rdata[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14811_ _14999_/A vssd1 vssd1 vccd1 vccd1 _14811_/X sky130_fd_sc_hd__buf_2
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15791_ _14996_/X _18905_/Q _15791_/S vssd1 vssd1 vccd1 vccd1 _15792_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11383__A _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17530_ _17530_/A vssd1 vssd1 vccd1 vccd1 _19626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14742_ _14742_/A vssd1 vssd1 vccd1 vccd1 _18588_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16929__A0 _16755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11954_ _11954_/A _11954_/B vssd1 vssd1 vccd1 vccd1 _11956_/A sky130_fd_sc_hd__nor2_2
X_10905_ _18588_/Q _19277_/Q _10905_/S vssd1 vssd1 vccd1 vccd1 _10906_/B sky130_fd_sc_hd__mux2_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17461_ _16844_/X _19596_/Q _17461_/S vssd1 vssd1 vccd1 vccd1 _17462_/A sky130_fd_sc_hd__mux2_1
X_14673_ _14673_/A vssd1 vssd1 vccd1 vccd1 _18207_/A sky130_fd_sc_hd__buf_4
XANTENNA__13207__A2 _12748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11885_ _17611_/B vssd1 vssd1 vccd1 vccd1 _11885_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16385__S _16391_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18166__A _18199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output108_A _13578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19200_ _19818_/CLK _19200_/D vssd1 vssd1 vccd1 vccd1 _19200_/Q sky130_fd_sc_hd__dfxtp_1
X_16412_ _16412_/A vssd1 vssd1 vccd1 vccd1 _19170_/D sky130_fd_sc_hd__clkbuf_1
X_13624_ _14057_/B _13623_/Y _13681_/S vssd1 vssd1 vccd1 vccd1 _13624_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12415__B1 _17693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10836_ _10836_/A _18854_/Q vssd1 vssd1 vccd1 vccd1 _10836_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17392_ _17448_/A vssd1 vssd1 vccd1 vccd1 _17461_/S sky130_fd_sc_hd__buf_8
XFILLER_158_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10426__C1 _09133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19131_ _19614_/CLK _19131_/D vssd1 vssd1 vccd1 vccd1 _19131_/Q sky130_fd_sc_hd__dfxtp_1
X_16343_ _16115_/X _19140_/Q _16351_/S vssd1 vssd1 vccd1 vccd1 _16344_/A sky130_fd_sc_hd__mux2_1
X_13555_ _13555_/A vssd1 vssd1 vccd1 vccd1 _18422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10767_ _09408_/A _10760_/Y _10762_/Y _10764_/Y _10766_/Y vssd1 vssd1 vccd1 vccd1
+ _10767_/X sky130_fd_sc_hd__o32a_1
XFILLER_41_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12506_ _13625_/A vssd1 vssd1 vccd1 vccd1 _13765_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_157_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16274_ _16274_/A vssd1 vssd1 vccd1 vccd1 _19109_/D sky130_fd_sc_hd__clkbuf_1
X_19062_ _19062_/CLK _19062_/D vssd1 vssd1 vccd1 vccd1 _19062_/Q sky130_fd_sc_hd__dfxtp_1
X_13486_ _18402_/Q _12634_/B _13486_/S vssd1 vssd1 vccd1 vccd1 _13487_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10698_ _10791_/A _10697_/X _09407_/A vssd1 vssd1 vccd1 vccd1 _10698_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_145_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18013_ _19789_/Q _18009_/B _18012_/Y vssd1 vssd1 vccd1 vccd1 _19789_/D sky130_fd_sc_hd__o21a_1
X_15225_ _15225_/A vssd1 vssd1 vccd1 vccd1 _18677_/D sky130_fd_sc_hd__clkbuf_1
X_12437_ _19689_/Q _11989_/X _12436_/Y _17711_/A vssd1 vssd1 vccd1 vccd1 _12437_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13391__A1 _18295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15156_ _15239_/S vssd1 vssd1 vccd1 vccd1 _15169_/S sky130_fd_sc_hd__buf_2
XFILLER_153_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12368_ _13388_/A _12393_/C vssd1 vssd1 vccd1 vccd1 _12368_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10824__S0 _11027_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12661__B _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14107_ _12008_/A _14111_/A vssd1 vssd1 vccd1 vccd1 _14107_/X sky130_fd_sc_hd__and2b_1
XFILLER_153_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11319_ _11471_/A _11376_/A _11551_/B _14547_/A vssd1 vssd1 vccd1 vccd1 _14274_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_4_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15087_ _18621_/Q _15086_/X _15087_/S vssd1 vssd1 vccd1 vccd1 _15088_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15132__A2 _13873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12299_ _13352_/A _12320_/C _17241_/S vssd1 vssd1 vccd1 vccd1 _12299_/X sky130_fd_sc_hd__a21o_1
XFILLER_141_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18915_ _19698_/CLK _18915_/D vssd1 vssd1 vccd1 vccd1 _18915_/Q sky130_fd_sc_hd__dfxtp_1
X_14038_ _13810_/A _13969_/X _13899_/A vssd1 vssd1 vccd1 vccd1 _14038_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_79_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15464__S _15470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10052__S1 _10029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18846_ _19624_/CLK _18846_/D vssd1 vssd1 vccd1 vccd1 _18846_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09993__S1 _09763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18777_ _19720_/CLK _18777_/D vssd1 vssd1 vccd1 vccd1 _18777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15989_ _15989_/A vssd1 vssd1 vccd1 vccd1 _18993_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17728_ _17728_/A _17728_/B vssd1 vssd1 vccd1 vccd1 _17728_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_40_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17659_ _17707_/A vssd1 vssd1 vccd1 vccd1 _17681_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09698__A _11157_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19329_ _19329_/CLK _19329_/D vssd1 vssd1 vccd1 vccd1 _19329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17896__A1 _19748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15639__S _15647_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09915_ _09163_/A _09913_/Y _09914_/Y _09770_/X vssd1 vssd1 vccd1 vccd1 _09915_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_98_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14882__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09846_ _09976_/A vssd1 vssd1 vccd1 vccd1 _09914_/A sky130_fd_sc_hd__clkbuf_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09777_ _18777_/Q _19006_/Q _18937_/Q _19235_/Q _09760_/X _09763_/X vssd1 vssd1 vccd1
+ vccd1 _09778_/B sky130_fd_sc_hd__mux4_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14634__A1 _18565_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16994__A _17062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11931__A _11984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _19661_/Q _12191_/A vssd1 vssd1 vccd1 vccd1 _11670_/X sky130_fd_sc_hd__or2_1
XFILLER_30_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10621_ _19509_/Q _19123_/Q _19573_/Q _18729_/Q _10353_/A _10366_/A vssd1 vssd1 vccd1
+ vccd1 _10622_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09401__A _10494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10547__A _10813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13340_ _18257_/Q _12651_/A _12752_/A _19782_/Q vssd1 vssd1 vccd1 vccd1 _13340_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17887__A1 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10552_ _09434_/A _10539_/X _10543_/X _10551_/X _10568_/A vssd1 vssd1 vccd1 vccd1
+ _10552_/X sky130_fd_sc_hd__a311o_2
XFILLER_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15898__A0 _14792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15549__S _15552_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13271_ _19482_/Q _13235_/X _13236_/X _18363_/Q _13270_/X vssd1 vssd1 vccd1 vccd1
+ _13273_/A sky130_fd_sc_hd__a221o_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10483_ _09275_/A _10473_/X _10482_/X _09282_/A _18437_/Q vssd1 vssd1 vccd1 vccd1
+ _11082_/B sky130_fd_sc_hd__a32o_4
XANTENNA__12762__A _14565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15010_ _15010_/A vssd1 vssd1 vccd1 vccd1 _15056_/S sky130_fd_sc_hd__buf_4
XFILLER_108_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12222_ _18371_/Q _18370_/Q _12222_/C vssd1 vssd1 vccd1 vccd1 _12272_/C sky130_fd_sc_hd__and3_1
XANTENNA__13373__A1 _19850_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10806__S0 _10932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10187__A1 _09867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input69_A io_irq_m3_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12153_ _11997_/A _12148_/Y _12151_/X _12152_/X vssd1 vssd1 vccd1 vccd1 _17890_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_118_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10282__S1 _11113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11104_ _09434_/X _11097_/X _11099_/X _11103_/X _09246_/A vssd1 vssd1 vccd1 vccd1
+ _11104_/X sky130_fd_sc_hd__a311o_2
XFILLER_96_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12084_ _12085_/A _13604_/A vssd1 vssd1 vccd1 vccd1 _12086_/A sky130_fd_sc_hd__and2_1
X_16961_ _16961_/A vssd1 vssd1 vccd1 vccd1 _19388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18700_ _19640_/CLK _18700_/D vssd1 vssd1 vccd1 vccd1 _18700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15912_ _15912_/A vssd1 vssd1 vccd1 vccd1 _18958_/D sky130_fd_sc_hd__clkbuf_1
X_11035_ _10821_/X _11026_/Y _11030_/Y _11034_/Y _09243_/A vssd1 vssd1 vccd1 vccd1
+ _11035_/X sky130_fd_sc_hd__o311a_2
X_19680_ _19680_/CLK _19680_/D vssd1 vssd1 vccd1 vccd1 _19680_/Q sky130_fd_sc_hd__dfxtp_1
X_16892_ _16892_/A vssd1 vssd1 vccd1 vccd1 _19358_/D sky130_fd_sc_hd__clkbuf_1
X_18631_ _19062_/CLK _18631_/D vssd1 vssd1 vccd1 vccd1 _18631_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_134_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15843_ _15865_/A vssd1 vssd1 vccd1 vccd1 _15852_/S sky130_fd_sc_hd__buf_4
XFILLER_40_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15822__A0 _14772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18562_ _19733_/CLK _18562_/D vssd1 vssd1 vccd1 vccd1 _18562_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _12997_/A _12993_/C vssd1 vssd1 vccd1 vccd1 _12986_/Y sky130_fd_sc_hd__nor2_1
X_15774_ _14908_/X _18897_/Q _15780_/S vssd1 vssd1 vccd1 vccd1 _15775_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ _17513_/A vssd1 vssd1 vccd1 vccd1 _19618_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ _11022_/X _13148_/B _14922_/S vssd1 vssd1 vccd1 vccd1 _14725_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ _11885_/X _11936_/Y _11801_/A vssd1 vssd1 vccd1 vccd1 _11937_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10111__A1 _10107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16378__A1 _15516_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18493_ _19468_/CLK _18493_/D vssd1 vssd1 vccd1 vccd1 _18493_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15313__A _15324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17444_ _16819_/X _19588_/Q _17446_/S vssd1 vssd1 vccd1 vccd1 _17445_/A sky130_fd_sc_hd__mux2_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14656_ _14696_/A vssd1 vssd1 vccd1 vccd1 _14677_/A sky130_fd_sc_hd__clkbuf_2
X_11868_ _11077_/A _18498_/Q _11948_/A vssd1 vssd1 vccd1 vccd1 _13617_/A sky130_fd_sc_hd__mux2_4
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12656__B _12656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10819_ _18757_/Q _18986_/Q _18917_/Q _19215_/Q _10905_/S _10739_/A vssd1 vssd1 vccd1
+ vccd1 _10820_/B sky130_fd_sc_hd__mux4_1
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13607_ _13607_/A vssd1 vssd1 vccd1 vccd1 _14126_/B sky130_fd_sc_hd__buf_2
X_17375_ _17375_/A vssd1 vssd1 vccd1 vccd1 _19557_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11799_ _11758_/X _11823_/B _18355_/Q vssd1 vssd1 vccd1 vccd1 _11799_/X sky130_fd_sc_hd__a21o_1
X_14587_ _14587_/A _14589_/B vssd1 vssd1 vccd1 vccd1 _14587_/X sky130_fd_sc_hd__or2_1
X_19114_ _19647_/CLK _19114_/D vssd1 vssd1 vccd1 vccd1 _19114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16326_ _16326_/A vssd1 vssd1 vccd1 vccd1 _19132_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13538_ _11552_/B _13536_/X _13537_/X _12555_/B vssd1 vssd1 vccd1 vccd1 _13539_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15889__A0 _14753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15459__S _15459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19045_ _19727_/CLK _19045_/D vssd1 vssd1 vccd1 vccd1 _19045_/Q sky130_fd_sc_hd__dfxtp_1
X_13469_ _18394_/Q _12713_/X _13475_/S vssd1 vssd1 vccd1 vccd1 _13470_/A sky130_fd_sc_hd__mux2_1
X_16257_ _16096_/X _19102_/Q _16257_/S vssd1 vssd1 vccd1 vccd1 _16258_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15208_ _18672_/Q _15207_/X _15217_/S vssd1 vssd1 vccd1 vccd1 _15209_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16188_ _16103_/X _19067_/Q _16194_/S vssd1 vssd1 vccd1 vccd1 _16189_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15139_ _15220_/A vssd1 vssd1 vccd1 vccd1 _15239_/S sky130_fd_sc_hd__buf_6
XFILLER_153_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14864__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09700_ _09700_/A vssd1 vssd1 vccd1 vccd1 _09701_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__09966__S1 _09936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09631_ _09631_/A vssd1 vssd1 vccd1 vccd1 _09632_/A sky130_fd_sc_hd__clkbuf_4
X_18829_ _19223_/CLK _18829_/D vssd1 vssd1 vccd1 vccd1 _18829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15813__A0 _14729_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15922__S _15924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10131__S _10131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ _09708_/A vssd1 vssd1 vccd1 vccd1 _09562_/X sky130_fd_sc_hd__buf_2
XFILLER_167_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16369__A1 _15503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09493_ _09493_/A vssd1 vssd1 vccd1 vccd1 _09493_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_3_0_0_clock_A clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15223__A _16725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15041__A1 _14744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09221__A _09856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17849__S _17849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15369__S _15373_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10169__A1 _10093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17584__S _17590_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15893__A _15950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11198__A _11199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09574__A3 _09573_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11926__A _11930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09957__S1 _09869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09829_ _09947_/A vssd1 vssd1 vccd1 vccd1 _09942_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ _18262_/Q _12840_/B _12840_/C vssd1 vssd1 vccd1 vccd1 _12841_/C sky130_fd_sc_hd__and3_1
XFILLER_73_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _13418_/S vssd1 vssd1 vccd1 vccd1 _13203_/A sky130_fd_sc_hd__buf_2
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11661__A _17221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11821_/A _12765_/A _11722_/C _11822_/B vssd1 vssd1 vccd1 vccd1 _11723_/C
+ sky130_fd_sc_hd__or4_1
X_14510_ _14510_/A vssd1 vssd1 vccd1 vccd1 _18523_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _15571_/A vssd1 vssd1 vccd1 vccd1 _15590_/S sky130_fd_sc_hd__clkbuf_16
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12476__B _12476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11653_ _11653_/A _11652_/X vssd1 vssd1 vccd1 vccd1 _11655_/A sky130_fd_sc_hd__or2b_2
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _18493_/Q _19731_/Q _14443_/S vssd1 vssd1 vccd1 vccd1 _14442_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10604_ _18594_/Q _19283_/Q _10604_/S vssd1 vssd1 vccd1 vccd1 _10604_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17160_ _17160_/A vssd1 vssd1 vccd1 vccd1 _19474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14372_ _18469_/Q vssd1 vssd1 vccd1 vccd1 _17662_/A sky130_fd_sc_hd__clkbuf_2
X_11584_ _11584_/A _11584_/B vssd1 vssd1 vccd1 vccd1 _13584_/D sky130_fd_sc_hd__and2_1
XFILLER_31_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16111_ _16111_/A vssd1 vssd1 vccd1 vccd1 _19037_/D sky130_fd_sc_hd__clkbuf_1
X_13323_ _12656_/B _13311_/X _13322_/X _13317_/X vssd1 vssd1 vccd1 vccd1 _18370_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10535_ _18827_/Q _19381_/Q _19543_/Q _18795_/Q _10560_/S _09634_/A vssd1 vssd1 vccd1
+ vccd1 _10535_/X sky130_fd_sc_hd__mux4_2
XFILLER_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13588__A _13720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17091_ _16781_/X _19446_/Q _17097_/S vssd1 vssd1 vccd1 vccd1 _17092_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13254_ _19866_/Q _12525_/X _12753_/X _19770_/Q vssd1 vssd1 vccd1 vccd1 _14824_/C
+ sky130_fd_sc_hd__a22o_2
X_16042_ _16752_/A vssd1 vssd1 vccd1 vccd1 _16042_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_8_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10466_ _18860_/Q _19318_/Q _10466_/S vssd1 vssd1 vccd1 vccd1 _10466_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09645__S0 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17494__S _17496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12205_ _14216_/A _12205_/B vssd1 vssd1 vccd1 vccd1 _12209_/A sky130_fd_sc_hd__xnor2_1
X_13185_ _13354_/A vssd1 vssd1 vccd1 vccd1 _13185_/X sky130_fd_sc_hd__clkbuf_2
X_10397_ _10438_/A _10396_/X _09315_/A vssd1 vssd1 vccd1 vccd1 _10397_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_123_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15099__A1 _18625_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19801_ _19804_/CLK _19801_/D vssd1 vssd1 vccd1 vccd1 _19801_/Q sky130_fd_sc_hd__dfxtp_1
X_12136_ _12137_/A _13596_/A vssd1 vssd1 vccd1 vccd1 _12138_/A sky130_fd_sc_hd__and2_1
XFILLER_150_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17993_ _17993_/A vssd1 vssd1 vccd1 vccd1 _17993_/X sky130_fd_sc_hd__buf_2
XFILLER_123_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19732_ _19732_/CLK _19732_/D vssd1 vssd1 vccd1 vccd1 _19732_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__11836__A _13761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12067_ _19741_/Q _12067_/B _19743_/Q _12067_/D vssd1 vssd1 vccd1 vccd1 _12092_/B
+ sky130_fd_sc_hd__and4_1
X_16944_ _16990_/S vssd1 vssd1 vccd1 vccd1 _16953_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__10740__A _10740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11018_ _18818_/Q _19372_/Q _19534_/Q _18786_/Q _10805_/A _10725_/A vssd1 vssd1 vccd1
+ vccd1 _11019_/B sky130_fd_sc_hd__mux4_1
X_19663_ _19682_/CLK _19663_/D vssd1 vssd1 vccd1 vccd1 _19663_/Q sky130_fd_sc_hd__dfxtp_2
X_16875_ _16875_/A vssd1 vssd1 vccd1 vccd1 _19350_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10332__A1 _19029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18614_ _19724_/CLK _18614_/D vssd1 vssd1 vccd1 vccd1 _18614_/Q sky130_fd_sc_hd__dfxtp_1
X_15826_ _14792_/X _18920_/Q _15830_/S vssd1 vssd1 vccd1 vccd1 _15827_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19594_ _19626_/CLK _19594_/D vssd1 vssd1 vccd1 vccd1 _19594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18545_ _19732_/CLK _18545_/D vssd1 vssd1 vccd1 vccd1 _18545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15757_ _15757_/A vssd1 vssd1 vccd1 vccd1 _18889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10886__S _10886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12667__A _12703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ _12972_/A _12972_/B _12922_/X vssd1 vssd1 vccd1 vccd1 _12969_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_33_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10096__B1 _09230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11571__A _19728_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15043__A _16731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14708_ _18458_/Q _14705_/X _14923_/S vssd1 vssd1 vccd1 vccd1 _14708_/X sky130_fd_sc_hd__mux2_2
XFILLER_127_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18476_ _18482_/CLK _18476_/D vssd1 vssd1 vccd1 vccd1 _18476_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15688_ _15734_/S vssd1 vssd1 vccd1 vccd1 _15697_/S sky130_fd_sc_hd__buf_2
XFILLER_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17427_ _16793_/X _19580_/Q _17435_/S vssd1 vssd1 vccd1 vccd1 _17428_/A sky130_fd_sc_hd__mux2_1
X_14639_ _14673_/A vssd1 vssd1 vccd1 vccd1 _14672_/A sky130_fd_sc_hd__buf_2
XANTENNA__16573__S _16573_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09976__A _09976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17358_ _17358_/A vssd1 vssd1 vccd1 vccd1 _19549_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15189__S _15201_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16309_ _16355_/S vssd1 vssd1 vccd1 vccd1 _16318_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__16523__A1 _15516_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10915__A _19693_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17289_ _19519_/Q _16699_/X _17291_/S vssd1 vssd1 vccd1 vccd1 _17290_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19028_ _19708_/CLK _19028_/D vssd1 vssd1 vccd1 vccd1 _19028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10246__S1 _10245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14837__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09216__A _10007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10323__B2 _18441_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15652__S _15658_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09614_ _11186_/S vssd1 vssd1 vccd1 vccd1 _09729_/S sky130_fd_sc_hd__buf_4
XFILLER_44_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ _18615_/Q _19304_/Q _09545_/S vssd1 vssd1 vccd1 vccd1 _09545_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09476_ _10579_/S vssd1 vssd1 vccd1 vccd1 _09522_/A sky130_fd_sc_hd__buf_2
XFILLER_12_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17579__S _17579_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4_0_clock_A clkbuf_4_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16514__A1 _15503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10320_ _11171_/A _10320_/B vssd1 vssd1 vccd1 vccd1 _10320_/X sky130_fd_sc_hd__or2_1
XFILLER_152_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_162_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10251_ _09402_/A _10234_/X _10250_/X vssd1 vssd1 vccd1 vccd1 _10251_/X sky130_fd_sc_hd__a21o_2
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09825__S _09874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10182_ _10182_/A _10182_/B vssd1 vssd1 vccd1 vccd1 _10182_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11656__A input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14990_ _14990_/A _15002_/C vssd1 vssd1 vccd1 vccd1 _14990_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13500__A1 _13364_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13941_ _13927_/A _13943_/B _13940_/X _13721_/X vssd1 vssd1 vccd1 vccd1 _13941_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_75_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15562__S _15568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17343__A _17389_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16660_ _16660_/A vssd1 vssd1 vccd1 vccd1 _19280_/D sky130_fd_sc_hd__clkbuf_1
X_13872_ _14328_/A _13851_/X _13869_/X _13871_/X vssd1 vssd1 vccd1 vccd1 _13872_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_90_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15611_ _15611_/A vssd1 vssd1 vccd1 vccd1 _18824_/D sky130_fd_sc_hd__clkbuf_1
X_12823_ _18257_/Q _18256_/Q _18255_/Q _12823_/D vssd1 vssd1 vccd1 vccd1 _12832_/D
+ sky130_fd_sc_hd__and4_1
X_16591_ _19251_/Q vssd1 vssd1 vccd1 vccd1 _16592_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_131_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12487__A _12487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11391__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18330_ _18330_/CLK _18330_/D vssd1 vssd1 vccd1 vccd1 _18330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_87_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15542_ _16797_/A vssd1 vssd1 vccd1 vccd1 _15542_/X sky130_fd_sc_hd__clkbuf_2
X_12754_ _18326_/Q _12663_/X _12753_/X _19783_/Q vssd1 vssd1 vccd1 vccd1 _12754_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15005__A1 _13363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ _19859_/CLK _18261_/D vssd1 vssd1 vccd1 vccd1 _18261_/Q sky130_fd_sc_hd__dfxtp_1
X_11705_ _12152_/B vssd1 vssd1 vccd1 vccd1 _11705_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15473_ _18778_/Q _15219_/X _15481_/S vssd1 vssd1 vccd1 vccd1 _15474_/A sky130_fd_sc_hd__mux2_1
X_12685_ _18622_/Q _12683_/Y _12684_/Y _12712_/A vssd1 vssd1 vccd1 vccd1 _13112_/A
+ sky130_fd_sc_hd__o22a_4
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _18447_/Q _13334_/X _17218_/S vssd1 vssd1 vccd1 vccd1 _17212_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09796__A _10153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14424_ _17765_/A _18519_/Q _14424_/S vssd1 vssd1 vccd1 vccd1 _14425_/A sky130_fd_sc_hd__mux2_1
X_11636_ _18576_/Q _14555_/A _11735_/S vssd1 vssd1 vccd1 vccd1 _11637_/C sky130_fd_sc_hd__mux2_1
X_18192_ _18249_/A _18192_/B _18196_/C vssd1 vssd1 vccd1 vccd1 _19851_/D sky130_fd_sc_hd__nor3_1
XFILLER_128_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17143_ _11022_/X _13149_/X _17143_/S vssd1 vssd1 vccd1 vccd1 _17143_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11567_ _12165_/S vssd1 vssd1 vccd1 vccd1 _12219_/S sky130_fd_sc_hd__clkbuf_2
X_14355_ _14384_/A vssd1 vssd1 vccd1 vccd1 _14367_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_128_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10476__S1 _10368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13306_ _13306_/A vssd1 vssd1 vccd1 vccd1 _13306_/X sky130_fd_sc_hd__clkbuf_2
X_10518_ _09529_/X _10513_/X _10517_/X _10589_/A vssd1 vssd1 vccd1 vccd1 _10518_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_157_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14286_ _14212_/A _14289_/B _13797_/X _14285_/X vssd1 vssd1 vccd1 vccd1 _14286_/X
+ sky130_fd_sc_hd__o211a_1
X_17074_ _17074_/A vssd1 vssd1 vccd1 vccd1 _19438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11498_ _18564_/Q _18562_/Q _11498_/C vssd1 vssd1 vccd1 vccd1 _11664_/D sky130_fd_sc_hd__or3_1
XFILLER_6_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09618__S0 _10131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13237_ _18276_/Q _13326_/B vssd1 vssd1 vccd1 vccd1 _13237_/X sky130_fd_sc_hd__and2_1
X_16025_ _15044_/X _19010_/Q _16027_/S vssd1 vssd1 vccd1 vccd1 _16026_/A sky130_fd_sc_hd__mux2_1
X_10449_ _10449_/A vssd1 vssd1 vccd1 vccd1 _10449_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10228__S1 _10390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13168_ _13139_/X _13165_/Y _13166_/X _13167_/X vssd1 vssd1 vccd1 vccd1 _18352_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10553__B2 _18436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ _14163_/A _12118_/Y _12119_/S vssd1 vssd1 vccd1 vccd1 _12119_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11566__A _11749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17976_ _19777_/Q _17979_/C _17950_/X vssd1 vssd1 vccd1 vccd1 _17976_/Y sky130_fd_sc_hd__a21oi_1
X_13099_ input68/X _13104_/B vssd1 vssd1 vccd1 vccd1 _13099_/X sky130_fd_sc_hd__or2_1
XFILLER_111_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15492__A1 _15487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19715_ _19715_/CLK _19715_/D vssd1 vssd1 vccd1 vccd1 _19715_/Q sky130_fd_sc_hd__dfxtp_1
X_16927_ _16752_/X _19373_/Q _16931_/S vssd1 vssd1 vccd1 vccd1 _16928_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19646_ _19712_/CLK _19646_/D vssd1 vssd1 vccd1 vccd1 _19646_/Q sky130_fd_sc_hd__dfxtp_1
X_16858_ _19343_/Q _16654_/X _16858_/S vssd1 vssd1 vccd1 vccd1 _16859_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15809_ _15865_/A vssd1 vssd1 vccd1 vccd1 _15878_/S sky130_fd_sc_hd__buf_8
X_19577_ _19609_/CLK _19577_/D vssd1 vssd1 vccd1 vccd1 _19577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16789_ _16789_/A vssd1 vssd1 vccd1 vccd1 _19320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09330_ _11180_/A vssd1 vssd1 vccd1 vccd1 _10140_/A sky130_fd_sc_hd__clkbuf_2
X_18528_ _18567_/CLK _18528_/D vssd1 vssd1 vccd1 vccd1 _18528_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11805__B2 _14578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10164__S0 _10200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09261_ _18420_/Q vssd1 vssd1 vccd1 vccd1 _16212_/C sky130_fd_sc_hd__clkbuf_2
X_18459_ _19693_/CLK _18459_/D vssd1 vssd1 vccd1 vccd1 _18459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09192_ _19693_/Q vssd1 vssd1 vccd1 vccd1 _10928_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09857__S0 _09163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10645__A _10764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10792__A1 _10634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15647__S _15647_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14286__A2 _14289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16478__S _16486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15382__S _15384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_109_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09528_ _19659_/Q _19076_/Q _19113_/Q _18719_/Q _10450_/S _09587_/A vssd1 vssd1 vccd1
+ vccd1 _09528_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _09459_/A vssd1 vssd1 vccd1 vccd1 _09459_/X sky130_fd_sc_hd__buf_2
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14726__S _14923_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17102__S _17108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12470_ _14545_/A _11313_/D _11664_/A vssd1 vssd1 vccd1 vccd1 _12471_/C sky130_fd_sc_hd__o21a_1
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11421_ _12519_/A _12520_/A _12747_/C vssd1 vssd1 vccd1 vccd1 _12516_/A sky130_fd_sc_hd__nor3_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14140_ _14297_/A _14140_/B vssd1 vssd1 vccd1 vccd1 _14140_/X sky130_fd_sc_hd__or2_1
X_11352_ _11375_/A _11640_/A vssd1 vssd1 vccd1 vccd1 _11476_/B sky130_fd_sc_hd__or2_2
XFILLER_126_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10783__B2 _12468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ _10309_/A vssd1 vssd1 vccd1 vccd1 _11166_/A sky130_fd_sc_hd__buf_2
X_14071_ _13881_/X _13886_/X _14085_/S vssd1 vssd1 vccd1 vccd1 _14071_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11283_ _11317_/A _11361_/A _11484_/A _11296_/C vssd1 vssd1 vccd1 vccd1 _13568_/B
+ sky130_fd_sc_hd__and4_1
X_13022_ _13024_/B _13024_/C _13021_/Y vssd1 vssd1 vccd1 vccd1 _18319_/D sky130_fd_sc_hd__o21a_1
XANTENNA_input51_A io_ibus_inst[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ _10219_/X _10222_/Y _10226_/Y _10229_/Y _10233_/Y vssd1 vssd1 vccd1 vccd1
+ _10234_/X sky130_fd_sc_hd__o32a_1
XFILLER_79_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17830_ _15203_/X _19716_/Q _17838_/S vssd1 vssd1 vccd1 vccd1 _17831_/A sky130_fd_sc_hd__mux2_1
X_10165_ _09996_/A _10164_/X _09215_/A vssd1 vssd1 vccd1 vccd1 _10165_/X sky130_fd_sc_hd__o21a_1
XFILLER_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17761_ _17765_/A _17765_/C vssd1 vssd1 vccd1 vccd1 _17761_/Y sky130_fd_sc_hd__xnor2_1
X_10096_ _10120_/A _10095_/X _09230_/A vssd1 vssd1 vccd1 vccd1 _10096_/X sky130_fd_sc_hd__o21a_1
X_14973_ _14969_/X _14971_/Y _14972_/Y vssd1 vssd1 vccd1 vccd1 _16712_/A sky130_fd_sc_hd__a21oi_4
XFILLER_47_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19500_ _19791_/CLK _19500_/D vssd1 vssd1 vccd1 vccd1 _19500_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15292__S _15300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16712_ _16712_/A vssd1 vssd1 vccd1 vccd1 _16712_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13924_ _13999_/S _13925_/B vssd1 vssd1 vccd1 vccd1 _13924_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17692_ _17701_/C _17692_/B vssd1 vssd1 vccd1 vccd1 _17692_/Y sky130_fd_sc_hd__nand2_1
X_19431_ _19724_/CLK _19431_/D vssd1 vssd1 vccd1 vccd1 _19431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16643_ _19275_/Q _16639_/X _16655_/S vssd1 vssd1 vccd1 vccd1 _16644_/A sky130_fd_sc_hd__mux2_1
X_13855_ _13810_/X _13854_/X _13819_/X vssd1 vssd1 vccd1 vccd1 _13855_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ _12991_/A vssd1 vssd1 vccd1 vccd1 _12851_/A sky130_fd_sc_hd__clkbuf_2
X_19362_ _19589_/CLK _19362_/D vssd1 vssd1 vccd1 vccd1 _19362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16574_ _16574_/A vssd1 vssd1 vccd1 vccd1 _19242_/D sky130_fd_sc_hd__clkbuf_1
X_10998_ _11026_/A _10997_/X _09223_/A vssd1 vssd1 vccd1 vccd1 _10998_/Y sky130_fd_sc_hd__o21ai_1
X_13786_ _13863_/A vssd1 vssd1 vccd1 vccd1 _14037_/A sky130_fd_sc_hd__clkbuf_2
X_18313_ _18330_/CLK _18313_/D vssd1 vssd1 vccd1 vccd1 _18313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15525_ _15525_/A vssd1 vssd1 vccd1 vccd1 _18795_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _12737_/A vssd1 vssd1 vccd1 vccd1 _12737_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19293_ _19616_/CLK _19293_/D vssd1 vssd1 vccd1 vccd1 _19293_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12945__A _18292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10697__S1 _10785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17012__S _17014_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18244_ _19869_/Q _18241_/B _18243_/Y vssd1 vssd1 vccd1 vccd1 _19869_/D sky130_fd_sc_hd__o21a_1
XFILLER_129_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15456_ _15456_/A vssd1 vssd1 vccd1 vccd1 _18770_/D sky130_fd_sc_hd__clkbuf_1
X_12668_ _13251_/A vssd1 vssd1 vccd1 vccd1 _12668_/X sky130_fd_sc_hd__buf_2
XFILLER_169_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14407_ _17737_/A _18513_/Q _14410_/S vssd1 vssd1 vccd1 vccd1 _14408_/A sky130_fd_sc_hd__mux2_1
X_18175_ _19845_/Q _19844_/Q _18175_/C vssd1 vssd1 vccd1 vccd1 _18177_/B sky130_fd_sc_hd__and3_1
XFILLER_128_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11619_ _11619_/A vssd1 vssd1 vccd1 vccd1 _11619_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15387_ _18741_/Q _15203_/X _15395_/S vssd1 vssd1 vccd1 vccd1 _15388_/A sky130_fd_sc_hd__mux2_1
X_12599_ _18339_/Q _12574_/X _12575_/X _12598_/X vssd1 vssd1 vccd1 vccd1 _18339_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_129_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17126_ _16832_/X _19462_/Q _17130_/S vssd1 vssd1 vccd1 vccd1 _17127_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14338_ _12450_/Y _13730_/X _14337_/X _15116_/A vssd1 vssd1 vccd1 vccd1 _14338_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17057_ _17057_/A vssd1 vssd1 vccd1 vccd1 _19431_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17248__A _17304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14269_ _13594_/X _13973_/Y _14268_/X _14097_/X vssd1 vssd1 vccd1 vccd1 _14269_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16152__A _16209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16008_ _14951_/X _19002_/Q _16016_/S vssd1 vssd1 vccd1 vccd1 _16009_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10621__S1 _10366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_191_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19640_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ _19770_/Q _17955_/C _17958_/Y vssd1 vssd1 vccd1 vccd1 _19770_/D sky130_fd_sc_hd__o21a_1
XFILLER_111_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_110_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__S0 _10277_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11743__B _11784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19629_ _19632_/CLK _19629_/D vssd1 vssd1 vccd1 vccd1 _19629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13016__A _13034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17711__A _17711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09313_ _09517_/A vssd1 vssd1 vccd1 vccd1 _09314_/A sky130_fd_sc_hd__buf_2
XFILLER_80_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10688__S1 _10670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09244_ _09244_/A vssd1 vssd1 vccd1 vccd1 _09245_/A sky130_fd_sc_hd__buf_2
X_09175_ _19693_/Q vssd1 vssd1 vccd1 vccd1 _10923_/A sky130_fd_sc_hd__inv_2
XANTENNA__12203__A1 _12491_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10214__A0 _19614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_144_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19630_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17158__A _17245_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_35_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11918__B _13622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16212__D _16212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10314__S _11156_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_159_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19599_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_163_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11190__A1 _09723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11934__A _19669_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11970_ _11970_/A vssd1 vssd1 vccd1 vccd1 _12106_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16001__S _16005_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10376__S0 _09448_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09404__A _09404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921_ _19503_/Q _19117_/Q _19567_/Q _18723_/Q _10919_/X _10920_/X vssd1 vssd1 vccd1
+ vccd1 _10922_/B sky130_fd_sc_hd__mux4_1
XFILLER_45_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13640_ _13776_/S vssd1 vssd1 vccd1 vccd1 _13743_/S sky130_fd_sc_hd__clkbuf_2
X_10852_ _18822_/Q _19376_/Q _19538_/Q _18790_/Q _10770_/S _09512_/A vssd1 vssd1 vccd1
+ vccd1 _10853_/B sky130_fd_sc_hd__mux4_2
XFILLER_72_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _10691_/X _12469_/A _11075_/A _12468_/A vssd1 vssd1 vccd1 vccd1 _11252_/A
+ sky130_fd_sc_hd__a22o_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _11643_/C _13571_/B _13571_/C _13571_/D vssd1 vssd1 vccd1 vccd1 _13572_/C
+ sky130_fd_sc_hd__and4b_1
XANTENNA__16237__A _16283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10679__S1 _09139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _15310_/A vssd1 vssd1 vccd1 vccd1 _18707_/D sky130_fd_sc_hd__clkbuf_1
X_12522_ _12602_/A vssd1 vssd1 vccd1 vccd1 _12522_/X sky130_fd_sc_hd__clkbuf_2
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16290_ _16039_/X _19116_/Q _16296_/S vssd1 vssd1 vccd1 vccd1 _16291_/A sky130_fd_sc_hd__mux2_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15241_ _15241_/A _15241_/B _15242_/C _15242_/D vssd1 vssd1 vccd1 vccd1 _15241_/X
+ sky130_fd_sc_hd__or4_4
X_12453_ _19690_/Q _13529_/B vssd1 vssd1 vccd1 vccd1 _12453_/X sky130_fd_sc_hd__or2_1
XFILLER_12_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16671__S _16671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11404_ _11404_/A vssd1 vssd1 vccd1 vccd1 _12747_/C sky130_fd_sc_hd__buf_2
X_15172_ _15239_/S vssd1 vssd1 vccd1 vccd1 _15185_/S sky130_fd_sc_hd__clkbuf_4
X_12384_ _12384_/A _12384_/B vssd1 vssd1 vccd1 vccd1 _12385_/B sky130_fd_sc_hd__nor2_2
XFILLER_138_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14123_ _13810_/X _13780_/X _13819_/X vssd1 vssd1 vccd1 vccd1 _14172_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__13596__A _13596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11335_ _11736_/B _14274_/A _13521_/B vssd1 vssd1 vccd1 vccd1 _13579_/A sky130_fd_sc_hd__or3b_1
XFILLER_67_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10851__S1 _10634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18931_ _19715_/CLK _18931_/D vssd1 vssd1 vccd1 vccd1 _18931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14054_ _14054_/A vssd1 vssd1 vccd1 vccd1 _14054_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11266_ _11266_/A _11266_/B _11266_/C _11266_/D vssd1 vssd1 vccd1 vccd1 _11266_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_134_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13005_ _17999_/A vssd1 vssd1 vccd1 vccd1 _13049_/A sky130_fd_sc_hd__clkbuf_2
X_10217_ _09215_/A _10210_/X _10212_/X _10216_/X _09248_/A vssd1 vssd1 vccd1 vccd1
+ _10217_/X sky130_fd_sc_hd__a311o_1
X_18862_ _19707_/CLK _18862_/D vssd1 vssd1 vccd1 vccd1 _18862_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12005__A _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11197_ _18454_/Q _09309_/A _09430_/A _11196_/X vssd1 vssd1 vccd1 vccd1 _12502_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_121_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17813_ _17813_/A vssd1 vssd1 vccd1 vccd1 _19708_/D sky130_fd_sc_hd__clkbuf_1
X_10148_ _18445_/Q vssd1 vssd1 vccd1 vccd1 _10148_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18793_ _19541_/CLK _18793_/D vssd1 vssd1 vccd1 vccd1 _18793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17744_ _17751_/C _17743_/Y _17711_/X vssd1 vssd1 vccd1 vccd1 _17744_/Y sky130_fd_sc_hd__a21oi_1
X_10079_ _19423_/Q _19199_/Q _19716_/Q _19167_/Q _10114_/S _09984_/A vssd1 vssd1 vccd1
+ vccd1 _10079_/X sky130_fd_sc_hd__mux4_1
X_14956_ _18479_/Q _14943_/X _14744_/X vssd1 vssd1 vccd1 vccd1 _14957_/B sky130_fd_sc_hd__o21ai_1
XFILLER_82_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13907_ _13795_/X _13903_/X _13904_/Y _13906_/X vssd1 vssd1 vccd1 vccd1 _13908_/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_36_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09314__A _09314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17675_ _17683_/C _17675_/B vssd1 vssd1 vccd1 vccd1 _17675_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14887_ _14887_/A _14887_/B vssd1 vssd1 vccd1 vccd1 _16689_/A sky130_fd_sc_hd__and2_2
XFILLER_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19414_ _19414_/CLK _19414_/D vssd1 vssd1 vccd1 vccd1 _19414_/Q sky130_fd_sc_hd__dfxtp_1
X_16626_ _16626_/A vssd1 vssd1 vccd1 vccd1 _19268_/D sky130_fd_sc_hd__clkbuf_1
X_13838_ _13838_/A vssd1 vssd1 vccd1 vccd1 _14135_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10119__S0 _10011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19345_ _19571_/CLK _19345_/D vssd1 vssd1 vccd1 vccd1 _19345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16557_ _16557_/A vssd1 vssd1 vccd1 vccd1 _19234_/D sky130_fd_sc_hd__clkbuf_1
X_13769_ _13767_/X _13768_/X _13769_/S vssd1 vssd1 vccd1 vccd1 _13769_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15508_ _18790_/Q _15506_/X _15520_/S vssd1 vssd1 vccd1 vccd1 _15509_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19276_ _19436_/CLK _19276_/D vssd1 vssd1 vccd1 vccd1 _19276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16488_ _16488_/A vssd1 vssd1 vccd1 vccd1 _16497_/S sky130_fd_sc_hd__buf_6
X_18227_ _19863_/Q _18223_/B _18226_/Y vssd1 vssd1 vccd1 vccd1 _19863_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_61_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19838_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15439_ _15485_/S vssd1 vssd1 vccd1 vccd1 _15448_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__10195__A _10196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18158_ _19840_/Q _18158_/B vssd1 vssd1 vccd1 vccd1 _18164_/C sky130_fd_sc_hd__and2_1
XFILLER_163_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17109_ _17109_/A vssd1 vssd1 vccd1 vccd1 _19454_/D sky130_fd_sc_hd__clkbuf_1
X_18089_ _18089_/A vssd1 vssd1 vccd1 vccd1 _18094_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10842__S1 _10785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16883__A0 _19354_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09931_ _09810_/X _09930_/X _09385_/A vssd1 vssd1 vccd1 vccd1 _09931_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_76_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19648_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_171_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09862_ _09237_/A _09859_/X _09861_/X _09231_/X vssd1 vssd1 vccd1 vccd1 _09862_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11172__A1 _11166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _09793_/A vssd1 vssd1 vccd1 vccd1 _09794_/A sky130_fd_sc_hd__buf_2
XFILLER_97_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15226__A _16728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12569__B _12715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15660__S _15662_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_14_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19580_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15610__A1 _15513_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13621__A0 _14074_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14177__A1 _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19715_/CLK sky130_fd_sc_hd__clkbuf_16
X_09227_ _09227_/A vssd1 vssd1 vccd1 vccd1 _09708_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__16491__S _16497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09158_ _11157_/S vssd1 vssd1 vccd1 vccd1 _11156_/S sky130_fd_sc_hd__buf_4
XFILLER_147_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09089_ _11339_/B vssd1 vssd1 vccd1 vccd1 _11376_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_163_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11120_ _19642_/Q _19059_/Q _19096_/Q _18702_/Q _10230_/X _10245_/X vssd1 vssd1 vccd1
+ vccd1 _11120_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11648__B _13650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15835__S _15841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11051_ _18849_/Q _19307_/Q _11051_/S vssd1 vssd1 vccd1 vccd1 _11052_/B sky130_fd_sc_hd__mux2_1
XFILLER_89_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11163__A1 _11166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15429__A1 _15155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ _09278_/X _09990_/X _10001_/X _09285_/X _18448_/Q vssd1 vssd1 vccd1 vccd1
+ _10003_/B sky130_fd_sc_hd__a32o_4
XFILLER_88_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14810_ _14810_/A vssd1 vssd1 vccd1 vccd1 _18594_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14101__A1 _18438_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15790_ _15790_/A vssd1 vssd1 vccd1 vccd1 _18904_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09134__A _09134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11383__B _13532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14741_ _14740_/X _18588_/Q _14762_/S vssd1 vssd1 vccd1 vccd1 _14742_/A sky130_fd_sc_hd__mux2_1
XANTENNA_input14_A io_dbus_rdata[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10123__C1 _09135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ _11953_/A _13620_/A vssd1 vssd1 vccd1 vccd1 _11954_/B sky130_fd_sc_hd__and2_1
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17460_ _17460_/A vssd1 vssd1 vccd1 vccd1 _19595_/D sky130_fd_sc_hd__clkbuf_1
X_10904_ _09427_/A _10893_/X _10902_/X _09625_/A _10903_/Y vssd1 vssd1 vccd1 vccd1
+ _12462_/A sky130_fd_sc_hd__o32a_4
XFILLER_72_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14672_ _14672_/A _15958_/B vssd1 vssd1 vccd1 vccd1 _18577_/D sky130_fd_sc_hd__nor2_1
X_11884_ _19667_/Q _12191_/A vssd1 vssd1 vccd1 vccd1 _11884_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15601__A1 _15500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16411_ _19170_/Q _15564_/X _16413_/S vssd1 vssd1 vccd1 vccd1 _16412_/A sky130_fd_sc_hd__mux2_1
X_13623_ _14216_/B vssd1 vssd1 vccd1 vccd1 _13623_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__12415__A1 _18379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17391_ _17391_/A _17391_/B vssd1 vssd1 vccd1 vccd1 _17448_/A sky130_fd_sc_hd__or2_2
X_10835_ _19312_/Q vssd1 vssd1 vccd1 vccd1 _10835_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19130_ _19612_/CLK _19130_/D vssd1 vssd1 vccd1 vccd1 _19130_/Q sky130_fd_sc_hd__dfxtp_1
X_16342_ _16342_/A vssd1 vssd1 vccd1 vccd1 _16351_/S sky130_fd_sc_hd__buf_6
XFILLER_13_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13554_ _13560_/A _13554_/B vssd1 vssd1 vccd1 vccd1 _13555_/A sky130_fd_sc_hd__and2_1
XFILLER_160_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10766_ _10762_/A _10765_/X _09408_/A vssd1 vssd1 vccd1 vccd1 _10766_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10977__A1 _10823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12505_ _12505_/A _12505_/B vssd1 vssd1 vccd1 vccd1 _12505_/Y sky130_fd_sc_hd__nor2_1
X_19061_ _19612_/CLK _19061_/D vssd1 vssd1 vccd1 vccd1 _19061_/Q sky130_fd_sc_hd__dfxtp_1
X_16273_ _16119_/X _19109_/Q _16279_/S vssd1 vssd1 vccd1 vccd1 _16274_/A sky130_fd_sc_hd__mux2_1
X_13485_ _13485_/A vssd1 vssd1 vccd1 vccd1 _18401_/D sky130_fd_sc_hd__clkbuf_1
X_10697_ _19636_/Q _19053_/Q _19090_/Q _18696_/Q _11050_/S _10785_/A vssd1 vssd1 vccd1
+ vccd1 _10697_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18012_ _18027_/A _18014_/B vssd1 vssd1 vccd1 vccd1 _18012_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15224_ _18677_/Q _15223_/X _15233_/S vssd1 vssd1 vccd1 vccd1 _15225_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12436_ _12294_/S _14319_/A _12435_/X vssd1 vssd1 vccd1 vccd1 _12436_/Y sky130_fd_sc_hd__o21bai_1
X_15155_ _16657_/A vssd1 vssd1 vccd1 vccd1 _15155_/X sky130_fd_sc_hd__buf_2
X_12367_ _13388_/A _12393_/C vssd1 vssd1 vccd1 vccd1 _12367_/X sky130_fd_sc_hd__or2_1
XANTENNA__10824__S1 _10813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10600__A_N _10601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14106_ _14019_/S _13850_/X _13706_/A vssd1 vssd1 vccd1 vccd1 _14106_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09309__A _09309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13679__A0 _12180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11318_ _11365_/A vssd1 vssd1 vccd1 vccd1 _14547_/A sky130_fd_sc_hd__clkbuf_2
X_12298_ _13352_/A _12320_/C vssd1 vssd1 vccd1 vccd1 _12298_/Y sky130_fd_sc_hd__nor2_1
X_15086_ _14555_/A _11070_/A _15092_/S vssd1 vssd1 vccd1 vccd1 _15086_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15745__S _15747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18914_ _19597_/CLK _18914_/D vssd1 vssd1 vccd1 vccd1 _18914_/Q sky130_fd_sc_hd__dfxtp_1
X_14037_ _14037_/A vssd1 vssd1 vccd1 vccd1 _14037_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11249_ _11249_/A vssd1 vssd1 vccd1 vccd1 _11249_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16430__A _16430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12351__A0 _09688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18845_ _19590_/CLK _18845_/D vssd1 vssd1 vccd1 vccd1 _18845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10362__C1 _09212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18776_ _19720_/CLK _18776_/D vssd1 vssd1 vccd1 vccd1 _18776_/Q sky130_fd_sc_hd__dfxtp_1
X_15988_ _14847_/X _18993_/Q _15994_/S vssd1 vssd1 vccd1 vccd1 _15989_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17727_ _17728_/A _17728_/B vssd1 vssd1 vccd1 vccd1 _17737_/C sky130_fd_sc_hd__or2_1
X_14939_ _16702_/A vssd1 vssd1 vccd1 vccd1 _16806_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_0_0_clock_A clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09979__A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17658_ _13259_/X _17657_/Y _17658_/S vssd1 vssd1 vccd1 vccd1 _17658_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16609_ _19260_/Q vssd1 vssd1 vccd1 vccd1 _16610_/A sky130_fd_sc_hd__clkbuf_1
X_17589_ _17589_/A vssd1 vssd1 vccd1 vccd1 _19652_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10918__A _19693_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19328_ _19620_/CLK _19328_/D vssd1 vssd1 vccd1 vccd1 _19328_/Q sky130_fd_sc_hd__dfxtp_1
X_19259_ _19613_/CLK _19259_/D vssd1 vssd1 vccd1 vccd1 _19259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10129__S _10129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11749__A _11749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09914_ _09914_/A _18872_/Q vssd1 vssd1 vccd1 vccd1 _09914_/Y sky130_fd_sc_hd__nor2_1
XFILLER_120_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14882__A2 _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _10115_/A _09844_/X _09788_/A vssd1 vssd1 vccd1 vccd1 _09845_/X sky130_fd_sc_hd__a21o_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A io_dbus_rdata[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09776_ _09861_/A _09764_/X _09767_/X _09775_/X vssd1 vssd1 vccd1 vccd1 _09776_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16486__S _16486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12645__A1 _19679_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10751__S0 _10669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10620_ _09210_/A _10603_/X _10607_/X _10619_/X _10568_/A vssd1 vssd1 vccd1 vccd1
+ _10620_/X sky130_fd_sc_hd__a311o_2
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10551_ _09549_/A _10544_/X _10550_/X _09459_/A vssd1 vssd1 vccd1 vccd1 _10551_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13270_ _18280_/Q _13270_/B vssd1 vssd1 vccd1 vccd1 _13270_/X sky130_fd_sc_hd__and2_1
X_10482_ _09212_/A _10475_/X _10477_/X _10481_/X _09246_/A vssd1 vssd1 vccd1 vccd1
+ _10482_/X sky130_fd_sc_hd__a311o_4
XANTENNA__11059__S1 _09480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12221_ _13322_/A _12222_/C _18371_/Q vssd1 vssd1 vccd1 vccd1 _12221_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11659__A _19730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10806__S1 _10713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12152_ _19746_/Q _12152_/B vssd1 vssd1 vccd1 vccd1 _12152_/X sky130_fd_sc_hd__or2_1
XFILLER_2_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09129__A _19695_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11103_ _09463_/A _11100_/X _11102_/X _09227_/A vssd1 vssd1 vccd1 vccd1 _11103_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15565__S _15568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16960_ _16800_/X _19388_/Q _16964_/S vssd1 vssd1 vccd1 vccd1 _16961_/A sky130_fd_sc_hd__mux2_1
X_12083_ _10299_/A _18506_/Q _12177_/A vssd1 vssd1 vccd1 vccd1 _13604_/A sky130_fd_sc_hd__mux2_4
XFILLER_151_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15911_ _14867_/X _18958_/Q _15913_/S vssd1 vssd1 vccd1 vccd1 _15912_/A sky130_fd_sc_hd__mux2_1
X_11034_ _11041_/A _11031_/X _11033_/X vssd1 vssd1 vccd1 vccd1 _11034_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16891_ _19358_/Q _16702_/X _16891_/S vssd1 vssd1 vccd1 vccd1 _16892_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10003__A_N _12493_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10344__C1 _09403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18630_ _19062_/CLK _18630_/D vssd1 vssd1 vccd1 vccd1 _18630_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_76_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15842_ _15842_/A vssd1 vssd1 vccd1 vccd1 _18927_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18561_ _18585_/CLK _18561_/D vssd1 vssd1 vccd1 vccd1 _18561_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15773_ _15773_/A vssd1 vssd1 vccd1 vccd1 _18896_/D sky130_fd_sc_hd__clkbuf_1
X_12985_ _12995_/D vssd1 vssd1 vccd1 vccd1 _12993_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16396__S _16402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14909__S _14941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_4_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ _19618_/Q _16709_/X _17518_/S vssd1 vssd1 vccd1 vccd1 _17513_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_157_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14724_ _14724_/A vssd1 vssd1 vccd1 vccd1 _18586_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ _18360_/Q _11936_/B vssd1 vssd1 vccd1 vccd1 _11936_/Y sky130_fd_sc_hd__xnor2_1
X_18492_ _18623_/CLK _18492_/D vssd1 vssd1 vccd1 vccd1 _18492_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10742__S0 _10669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17443_ _17443_/A vssd1 vssd1 vccd1 vccd1 _19587_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14655_ _14655_/A vssd1 vssd1 vccd1 vccd1 _18571_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _14026_/A _11867_/B vssd1 vssd1 vccd1 vccd1 _11870_/A sky130_fd_sc_hd__xor2_1
X_13606_ _14138_/B _14155_/B _13685_/S vssd1 vssd1 vccd1 vccd1 _13606_/X sky130_fd_sc_hd__mux2_1
X_17374_ _16822_/X _19557_/Q _17374_/S vssd1 vssd1 vccd1 vccd1 _17375_/A sky130_fd_sc_hd__mux2_1
X_10818_ _19407_/Q _19183_/Q _19700_/Q _19151_/Q _10982_/S _10969_/A vssd1 vssd1 vccd1
+ vccd1 _10818_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14586_ _18551_/Q _14577_/X _14584_/X _14585_/X vssd1 vssd1 vccd1 vccd1 _18551_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11798_ _18355_/Q _11823_/B vssd1 vssd1 vccd1 vccd1 _11798_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19113_ _19659_/CLK _19113_/D vssd1 vssd1 vccd1 vccd1 _19113_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11630__D_N _11624_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16325_ _16090_/X _19132_/Q _16329_/S vssd1 vssd1 vccd1 vccd1 _16326_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13537_ _13537_/A vssd1 vssd1 vccd1 vccd1 _13537_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12953__A _12983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10749_ _19635_/Q _19052_/Q _19089_/Q _18695_/Q _10669_/A _10670_/X vssd1 vssd1 vccd1
+ vccd1 _10750_/B sky130_fd_sc_hd__mux4_1
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19044_ _19713_/CLK _19044_/D vssd1 vssd1 vccd1 vccd1 _19044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16256_ _16256_/A vssd1 vssd1 vccd1 vccd1 _19101_/D sky130_fd_sc_hd__clkbuf_1
X_13468_ _13468_/A vssd1 vssd1 vccd1 vccd1 _18393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15207_ _16709_/A vssd1 vssd1 vccd1 vccd1 _15207_/X sky130_fd_sc_hd__clkbuf_2
X_12419_ _12419_/A _12419_/B vssd1 vssd1 vccd1 vccd1 _14324_/A sky130_fd_sc_hd__nand2_4
XFILLER_173_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16187_ _16187_/A vssd1 vssd1 vccd1 vccd1 _19066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13399_ _12577_/X _13390_/Y _13398_/X _12596_/X _18647_/Q vssd1 vssd1 vccd1 vccd1
+ _13399_/X sky130_fd_sc_hd__a32o_4
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15138_ _17463_/A _16847_/B vssd1 vssd1 vccd1 vccd1 _15220_/A sky130_fd_sc_hd__nor2_2
XFILLER_126_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15475__S _15481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14313__A1 _14310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15069_ _18489_/Q _15069_/B vssd1 vssd1 vccd1 vccd1 _15069_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14864__A2 _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09630_ _10560_/S vssd1 vssd1 vccd1 vccd1 _09631_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18828_ _19543_/CLK _18828_/D vssd1 vssd1 vccd1 vccd1 _18828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09561_ _09649_/A _09561_/B vssd1 vssd1 vccd1 vccd1 _09561_/X sky130_fd_sc_hd__or2_1
X_18759_ _19442_/CLK _18759_/D vssd1 vssd1 vccd1 vccd1 _18759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09492_ _18879_/Q _19337_/Q _10511_/S vssd1 vssd1 vccd1 vccd1 _09493_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17566__A1 _16787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11751__B _11751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11470__C _14431_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_4_0_clock_A clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11198__B _12502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13107__A2 _12731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09731__A1 _10132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09828_ _10042_/A vssd1 vssd1 vccd1 vccd1 _09947_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14607__A2 _13106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10972__S0 _10919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09759_ _10076_/S vssd1 vssd1 vccd1 vccd1 _10075_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15414__A _16992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13291__A1 _19838_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12770_ _12765_/A _13108_/A _13115_/A _18374_/Q _12769_/X vssd1 vssd1 vccd1 vccd1
+ _12770_/X sky130_fd_sc_hd__a221o_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09412__A _09412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _11721_/A _11444_/X vssd1 vssd1 vccd1 vccd1 _11721_/X sky130_fd_sc_hd__or2b_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14440_/A vssd1 vssd1 vccd1 vccd1 _18492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11652_ _11652_/A _13665_/A vssd1 vssd1 vccd1 vccd1 _11652_/X sky130_fd_sc_hd__or2_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10603_ _10622_/A _10603_/B vssd1 vssd1 vccd1 vccd1 _10603_/X sky130_fd_sc_hd__or2_1
XFILLER_128_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14371_ _14371_/A vssd1 vssd1 vccd1 vccd1 _18468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11583_ _13583_/B _11585_/D vssd1 vssd1 vccd1 vccd1 _11644_/A sky130_fd_sc_hd__nor2_1
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16110_ _16109_/X _19037_/Q _16113_/S vssd1 vssd1 vccd1 vccd1 _16111_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13322_ _13322_/A _13352_/B vssd1 vssd1 vccd1 vccd1 _13322_/X sky130_fd_sc_hd__or2_1
X_17090_ _17090_/A vssd1 vssd1 vccd1 vccd1 _19445_/D sky130_fd_sc_hd__clkbuf_1
X_10534_ _10566_/A _10534_/B vssd1 vssd1 vccd1 vccd1 _10534_/X sky130_fd_sc_hd__or2_1
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16041_ _16041_/A vssd1 vssd1 vccd1 vccd1 _19015_/D sky130_fd_sc_hd__clkbuf_1
X_13253_ _13253_/A _13253_/B vssd1 vssd1 vccd1 vccd1 _14824_/B sky130_fd_sc_hd__or2_1
X_10465_ _18597_/Q _19286_/Q _10465_/S vssd1 vssd1 vccd1 vccd1 _10465_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12204_ _12057_/A _14203_/A _12176_/B vssd1 vssd1 vccd1 vccd1 _12205_/B sky130_fd_sc_hd__a21oi_1
XFILLER_136_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13184_ _13139_/X _13182_/X _13183_/X _13167_/X vssd1 vssd1 vccd1 vccd1 _18354_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10396_ _19417_/Q _19193_/Q _19710_/Q _19161_/Q _09673_/S _09602_/A vssd1 vssd1 vccd1
+ vccd1 _10396_/X sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_83_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15099__A2 _13566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19800_ _19804_/CLK _19800_/D vssd1 vssd1 vccd1 vccd1 _19800_/Q sky130_fd_sc_hd__dfxtp_1
X_12135_ _10196_/A _18508_/Q _12328_/A vssd1 vssd1 vccd1 vccd1 _13596_/A sky130_fd_sc_hd__mux2_4
X_17992_ _19782_/Q _17990_/B _17991_/Y vssd1 vssd1 vccd1 vccd1 _19782_/D sky130_fd_sc_hd__o21a_1
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12306__A0 _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19731_ _19732_/CLK _19731_/D vssd1 vssd1 vccd1 vccd1 _19731_/Q sky130_fd_sc_hd__dfxtp_4
X_16943_ _16943_/A vssd1 vssd1 vccd1 vccd1 _19380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12066_ _12066_/A _12066_/B vssd1 vssd1 vccd1 vccd1 _12066_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__14212__B _14216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11017_ _19598_/Q _19436_/Q _18882_/Q _18652_/Q _10710_/A _09480_/A vssd1 vssd1 vccd1
+ vccd1 _11017_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19662_ _19689_/CLK _19662_/D vssd1 vssd1 vccd1 vccd1 _19662_/Q sky130_fd_sc_hd__dfxtp_2
X_16874_ _19350_/Q _16677_/X _16880_/S vssd1 vssd1 vccd1 vccd1 _16875_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15825_ _15825_/A vssd1 vssd1 vccd1 vccd1 _18919_/D sky130_fd_sc_hd__clkbuf_1
X_18613_ _19723_/CLK _18613_/D vssd1 vssd1 vccd1 vccd1 _18613_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12609__A1 _19487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19593_ _19657_/CLK _19593_/D vssd1 vssd1 vccd1 vccd1 _19593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12948__A _17895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15324__A _15324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18544_ _19732_/CLK _18544_/D vssd1 vssd1 vccd1 vccd1 _18544_/Q sky130_fd_sc_hd__dfxtp_1
X_15756_ _14808_/X _18889_/Q _15758_/S vssd1 vssd1 vccd1 vccd1 _15757_/A sky130_fd_sc_hd__mux2_1
X_12968_ _18304_/Q vssd1 vssd1 vccd1 vccd1 _12972_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10715__S0 _10706_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16139__B _16920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14707_ _14825_/A vssd1 vssd1 vccd1 vccd1 _14923_/S sky130_fd_sc_hd__buf_2
XFILLER_33_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11919_ _11919_/A _11919_/B vssd1 vssd1 vccd1 vccd1 _11920_/A sky130_fd_sc_hd__nand2_1
X_18475_ _18482_/CLK _18475_/D vssd1 vssd1 vccd1 vccd1 _18475_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15687_ _15687_/A vssd1 vssd1 vccd1 vccd1 _18858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12899_ _18279_/Q vssd1 vssd1 vccd1 vccd1 _12910_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _17448_/A vssd1 vssd1 vccd1 vccd1 _17435_/S sky130_fd_sc_hd__buf_4
X_14638_ _14638_/A _14638_/B vssd1 vssd1 vccd1 vccd1 _18566_/D sky130_fd_sc_hd__nor2_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17357_ _16797_/X _19549_/Q _17363_/S vssd1 vssd1 vccd1 vccd1 _17358_/A sky130_fd_sc_hd__mux2_1
X_14569_ _12533_/B _14564_/X _14568_/X _14560_/X vssd1 vssd1 vccd1 vccd1 _18544_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12683__A _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16308_ _16308_/A vssd1 vssd1 vccd1 vccd1 _19124_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17288_ _17288_/A vssd1 vssd1 vccd1 vccd1 _19518_/D sky130_fd_sc_hd__clkbuf_1
X_19027_ _19610_/CLK _19027_/D vssd1 vssd1 vccd1 vccd1 _19027_/Q sky130_fd_sc_hd__dfxtp_1
X_16239_ _16239_/A vssd1 vssd1 vccd1 vccd1 _19093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11_0_clock_A clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15933__S _15935_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10323__A2 _10311_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09613_ _09661_/A vssd1 vssd1 vccd1 vccd1 _11178_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_141_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ _09793_/A vssd1 vssd1 vccd1 vccd1 _09545_/S sky130_fd_sc_hd__buf_4
XFILLER_24_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09475_ _10591_/A vssd1 vssd1 vccd1 vccd1 _10392_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15970__A0 _14753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13328__A2 _12668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17595__S _17601_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_8_0_clock_A clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10250_ _09681_/X _10236_/Y _10244_/X _10249_/Y _09393_/A vssd1 vssd1 vccd1 vccd1
+ _10250_/X sky130_fd_sc_hd__o311a_1
XFILLER_105_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10181_ _19261_/Q _19032_/Q _18963_/Q _19357_/Q _10131_/S _09610_/X vssd1 vssd1 vccd1
+ vccd1 _10182_/B sky130_fd_sc_hd__mux4_1
XFILLER_59_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09407__A _09407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12839__A1 _12840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13940_ _13937_/X _13936_/B _14088_/A _13939_/X vssd1 vssd1 vccd1 vccd1 _13940_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10945__S0 _10706_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13871_ _14115_/A vssd1 vssd1 vccd1 vccd1 _13871_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12768__A _13154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15610_ _18824_/Q _15513_/X _15614_/S vssd1 vssd1 vccd1 vccd1 _15611_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12822_ _12851_/A _12822_/B _12822_/C vssd1 vssd1 vccd1 vccd1 _18256_/D sky130_fd_sc_hd__nor3_1
XFILLER_28_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13264__A1 _12713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16590_ _16590_/A vssd1 vssd1 vccd1 vccd1 _19250_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14461__A0 _18502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10078__A1 _09783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09142__A _09142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_opt_3_0_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15541_ _15541_/A vssd1 vssd1 vccd1 vccd1 _18800_/D sky130_fd_sc_hd__clkbuf_1
X_12753_ _12753_/A vssd1 vssd1 vccd1 vccd1 _12753_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _19859_/CLK _18260_/D vssd1 vssd1 vccd1 vccd1 _18260_/Q sky130_fd_sc_hd__dfxtp_1
X_11704_ _11746_/B _11704_/B vssd1 vssd1 vccd1 vccd1 _11704_/Y sky130_fd_sc_hd__nor2_8
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15472_ _15472_/A vssd1 vssd1 vccd1 vccd1 _15481_/S sky130_fd_sc_hd__buf_6
X_12684_ _12766_/A _18622_/Q _12600_/A vssd1 vssd1 vccd1 vccd1 _12684_/Y sky130_fd_sc_hd__a21boi_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17211_/A vssd1 vssd1 vccd1 vccd1 _19489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _18487_/Q vssd1 vssd1 vccd1 vccd1 _17765_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13599__A _13643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18191_ _19851_/Q _19850_/Q _18191_/C vssd1 vssd1 vccd1 vccd1 _18196_/C sky130_fd_sc_hd__and3_1
X_11635_ _18571_/Q vssd1 vssd1 vccd1 vccd1 _14555_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11122__S0 _09583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17142_ _17142_/A vssd1 vssd1 vccd1 vccd1 _19469_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12775__B1 _12748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09432__A1_N _18457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14354_ _18463_/Q vssd1 vssd1 vccd1 vccd1 _17632_/A sky130_fd_sc_hd__buf_2
XFILLER_155_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11566_ _11749_/A vssd1 vssd1 vccd1 vccd1 _12165_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_10_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13305_ _18634_/Q _13305_/B vssd1 vssd1 vccd1 vccd1 _13305_/X sky130_fd_sc_hd__or2_1
XANTENNA__10250__A1 _09681_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17073_ _16755_/X _19438_/Q _17075_/S vssd1 vssd1 vccd1 vccd1 _17074_/A sky130_fd_sc_hd__mux2_1
X_10517_ _09679_/A _10514_/X _10516_/X _09314_/A vssd1 vssd1 vccd1 vccd1 _10517_/X
+ sky130_fd_sc_hd__o211a_1
X_14285_ _14285_/A _14289_/A vssd1 vssd1 vccd1 vccd1 _14285_/X sky130_fd_sc_hd__or2_1
XFILLER_156_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11497_ _11497_/A _18565_/Q _18563_/Q vssd1 vssd1 vccd1 vccd1 _11498_/C sky130_fd_sc_hd__or3_1
XFILLER_171_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09618__S1 _09610_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16024_ _16024_/A vssd1 vssd1 vccd1 vccd1 _19009_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13236_ _13236_/A vssd1 vssd1 vccd1 vccd1 _13236_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10448_ _18861_/Q _19319_/Q _10486_/S vssd1 vssd1 vccd1 vccd1 _10449_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10002__B2 _18448_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11847__A _14431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ _17781_/A vssd1 vssd1 vccd1 vccd1 _13167_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14223__A _14227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10379_ _10379_/A _10379_/B vssd1 vssd1 vccd1 vccd1 _10379_/X sky130_fd_sc_hd__or2_1
XFILLER_112_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10553__A2 _10537_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12118_ _19745_/Q _12144_/C vssd1 vssd1 vccd1 vccd1 _12118_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09317__A _09317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13098_ _18343_/Q _12731_/X _13094_/X _14612_/A vssd1 vssd1 vccd1 vccd1 _18343_/D
+ sky130_fd_sc_hd__o211a_1
X_17975_ _19776_/Q _17973_/B _17974_/Y vssd1 vssd1 vccd1 vccd1 _19776_/D sky130_fd_sc_hd__o21a_1
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17218__A0 _18449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19714_ _19714_/CLK _19714_/D vssd1 vssd1 vccd1 vccd1 _19714_/Q sky130_fd_sc_hd__dfxtp_1
X_12049_ _18364_/Q vssd1 vssd1 vccd1 vccd1 _13295_/A sky130_fd_sc_hd__clkbuf_2
X_16926_ _16926_/A vssd1 vssd1 vccd1 vccd1 _19372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17769__A1 _19689_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10936__S0 _10886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19645_ _19645_/CLK _19645_/D vssd1 vssd1 vccd1 vccd1 _19645_/Q sky130_fd_sc_hd__dfxtp_1
X_16857_ _16857_/A vssd1 vssd1 vccd1 vccd1 _19342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15054__A _16734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15808_ _17391_/A _16503_/B vssd1 vssd1 vccd1 vccd1 _15865_/A sky130_fd_sc_hd__or2_2
XFILLER_80_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19576_ _19608_/CLK _19576_/D vssd1 vssd1 vccd1 vccd1 _19576_/Q sky130_fd_sc_hd__dfxtp_1
X_16788_ _16787_/X _19320_/Q _16791_/S vssd1 vssd1 vccd1 vccd1 _16789_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18527_ _18564_/CLK _18527_/D vssd1 vssd1 vccd1 vccd1 _18527_/Q sky130_fd_sc_hd__dfxtp_1
X_15739_ _14714_/X _18881_/Q _15747_/S vssd1 vssd1 vccd1 vccd1 _15740_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14893__A _14893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10164__S1 _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09260_ _18572_/Q _14716_/A vssd1 vssd1 vccd1 vccd1 _09260_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18458_ _19693_/CLK _18458_/D vssd1 vssd1 vccd1 vccd1 _18458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09191_ _19274_/Q _19045_/Q _18976_/Q _19370_/Q _09190_/X _09149_/A vssd1 vssd1 vccd1
+ vccd1 _09191_/X sky130_fd_sc_hd__mux4_1
X_17409_ _16768_/X _19572_/Q _17413_/S vssd1 vssd1 vccd1 vccd1 _17410_/A sky130_fd_sc_hd__mux2_1
X_18389_ _19689_/CLK _18389_/D vssd1 vssd1 vccd1 vccd1 _18389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11757__A _12715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15229__A _16731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11492__A _14589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_31_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09527_ _10496_/A _09527_/B vssd1 vssd1 vccd1 vccd1 _09527_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12454__C1 _17711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09897__A _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09458_ _10574_/A _09458_/B vssd1 vssd1 vccd1 vccd1 _09458_/X sky130_fd_sc_hd__or2_1
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10836__A _10836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09389_ _18981_/Q vssd1 vssd1 vccd1 vccd1 _09390_/A sky130_fd_sc_hd__inv_2
XFILLER_40_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14308__A _14310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11420_ _12670_/C _12540_/B _12563_/A _12585_/A _12603_/A vssd1 vssd1 vccd1 vccd1
+ _11427_/B sky130_fd_sc_hd__a2111o_1
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09622__B1 _09621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10555__B _12476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11351_ _11356_/A vssd1 vssd1 vccd1 vccd1 _11640_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_138_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10783__A2 _12469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10302_ _10313_/A _10302_/B vssd1 vssd1 vccd1 vccd1 _10302_/X sky130_fd_sc_hd__or2_1
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14070_ _14070_/A vssd1 vssd1 vccd1 vccd1 _14070_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11282_ _11282_/A vssd1 vssd1 vccd1 vccd1 _14545_/A sky130_fd_sc_hd__clkbuf_2
X_13021_ _13024_/B _13024_/C _13011_/X vssd1 vssd1 vccd1 vccd1 _13021_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10233_ _10226_/A _10232_/X _10219_/X vssd1 vssd1 vccd1 vccd1 _10233_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_117_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input44_A io_ibus_inst[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10164_ _19647_/Q _19064_/Q _19101_/Q _18707_/Q _10200_/S _09979_/A vssd1 vssd1 vccd1
+ vccd1 _10164_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17354__A _17376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17760_ _19687_/Q _17708_/A _17758_/Y _17759_/X vssd1 vssd1 vccd1 vccd1 _19687_/D
+ sky130_fd_sc_hd__o22a_1
X_10095_ _19617_/Q _19455_/Q _18901_/Q _18671_/Q _10094_/X _09769_/A vssd1 vssd1 vccd1
+ vccd1 _10095_/X sky130_fd_sc_hd__mux4_1
X_14972_ input15/X _14901_/X _14904_/X vssd1 vssd1 vccd1 vccd1 _14972_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16711_ _16711_/A vssd1 vssd1 vccd1 vccd1 _19296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13923_ _13942_/A vssd1 vssd1 vccd1 vccd1 _14078_/A sky130_fd_sc_hd__buf_2
XFILLER_47_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17691_ _18474_/Q _17691_/B vssd1 vssd1 vccd1 vccd1 _17692_/B sky130_fd_sc_hd__nand2_1
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12498__A _12505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16642_ _16741_/S vssd1 vssd1 vccd1 vccd1 _16655_/S sky130_fd_sc_hd__buf_2
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19430_ _19624_/CLK _19430_/D vssd1 vssd1 vccd1 vccd1 _19430_/Q sky130_fd_sc_hd__dfxtp_1
X_13854_ _13750_/X _13853_/X _13816_/X vssd1 vssd1 vccd1 vccd1 _13854_/X sky130_fd_sc_hd__o21a_1
XFILLER_35_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12805_ _13042_/A vssd1 vssd1 vccd1 vccd1 _12991_/A sky130_fd_sc_hd__buf_2
XFILLER_62_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09536__S0 _11157_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13106__B _13106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19361_ _19833_/CLK _19361_/D vssd1 vssd1 vccd1 vccd1 _19361_/Q sky130_fd_sc_hd__dfxtp_1
X_16573_ _19242_/Q _15589_/X _16573_/S vssd1 vssd1 vccd1 vccd1 _16574_/A sky130_fd_sc_hd__mux2_1
X_13785_ _13785_/A _13922_/B vssd1 vssd1 vccd1 vccd1 _13863_/A sky130_fd_sc_hd__or2_1
XFILLER_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10997_ _19598_/Q _19436_/Q _18882_/Q _18652_/Q _10663_/A _10364_/A vssd1 vssd1 vccd1
+ vccd1 _10997_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12010__B _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18312_ _19795_/CLK _18312_/D vssd1 vssd1 vccd1 vccd1 _18312_/Q sky130_fd_sc_hd__dfxtp_1
X_15524_ _18795_/Q _15522_/X _15536_/S vssd1 vssd1 vccd1 vccd1 _15525_/A sky130_fd_sc_hd__mux2_1
X_12736_ _12736_/A vssd1 vssd1 vccd1 vccd1 _12736_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19292_ _19613_/CLK _19292_/D vssd1 vssd1 vccd1 vccd1 _19292_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _18250_/A _18247_/C vssd1 vssd1 vccd1 vccd1 _18243_/Y sky130_fd_sc_hd__nor2_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15455_ _18770_/Q _15194_/X _15459_/S vssd1 vssd1 vccd1 vccd1 _15456_/A sky130_fd_sc_hd__mux2_1
X_12667_ _12703_/A vssd1 vssd1 vccd1 vccd1 _13251_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13122__A _13171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14406_ _18481_/Q vssd1 vssd1 vccd1 vccd1 _17737_/A sky130_fd_sc_hd__clkbuf_2
X_18174_ _19844_/Q _18175_/C _19845_/Q vssd1 vssd1 vccd1 vccd1 _18176_/B sky130_fd_sc_hd__a21oi_1
X_11618_ _11618_/A _11618_/B _11688_/C vssd1 vssd1 vccd1 vccd1 _11622_/B sky130_fd_sc_hd__and3_1
X_15386_ _15397_/A vssd1 vssd1 vccd1 vccd1 _15395_/S sky130_fd_sc_hd__buf_4
X_12598_ _12575_/X _12598_/B vssd1 vssd1 vccd1 vccd1 _12598_/X sky130_fd_sc_hd__and2b_1
X_17125_ _17125_/A vssd1 vssd1 vccd1 vccd1 _19461_/D sky130_fd_sc_hd__clkbuf_1
X_14337_ _13594_/X _13706_/Y _14097_/A _14336_/X vssd1 vssd1 vccd1 vccd1 _14337_/X
+ sky130_fd_sc_hd__o211a_1
X_11549_ _11549_/A vssd1 vssd1 vccd1 vccd1 _11552_/A sky130_fd_sc_hd__inv_2
XFILLER_143_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16433__A _16501_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17056_ _19431_/Q _16731_/X _17058_/S vssd1 vssd1 vccd1 vccd1 _17057_/A sky130_fd_sc_hd__mux2_1
X_14268_ _13971_/X _13970_/X _14267_/X vssd1 vssd1 vccd1 vccd1 _14268_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13173__B1 _12671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16007_ _16018_/A vssd1 vssd1 vccd1 vccd1 _16016_/S sky130_fd_sc_hd__buf_4
XFILLER_98_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13219_ _19832_/Q vssd1 vssd1 vccd1 vccd1 _18140_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_125_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _14203_/A _14203_/B vssd1 vssd1 vccd1 vccd1 _14199_/Y sky130_fd_sc_hd__nand2_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14888__A _16689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15483__S _15485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17958_ _17991_/A _17963_/C vssd1 vssd1 vccd1 vccd1 _17958_/Y sky130_fd_sc_hd__nor2_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16909_ _19366_/Q _16728_/X _16913_/S vssd1 vssd1 vccd1 vccd1 _16910_/A sky130_fd_sc_hd__mux2_1
X_17889_ _17889_/A vssd1 vssd1 vccd1 vccd1 _19745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19628_ _19628_/CLK _19628_/D vssd1 vssd1 vccd1 vccd1 _19628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19559_ _19559_/CLK _19559_/D vssd1 vssd1 vccd1 vccd1 _19559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09312_ _10793_/A vssd1 vssd1 vccd1 vccd1 _09517_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09510__A _09522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ _09243_/A vssd1 vssd1 vccd1 vccd1 _09244_/A sky130_fd_sc_hd__buf_2
XFILLER_166_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09174_ _18880_/Q _19338_/Q _09190_/A vssd1 vssd1 vccd1 vccd1 _09174_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15658__S _15658_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11487__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16489__S _16497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15393__S _15395_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13467__A1 _13259_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14310__B _14310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10376__S1 _09554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17902__A _19752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ _10960_/A vssd1 vssd1 vccd1 vccd1 _10920_/X sky130_fd_sc_hd__buf_4
XANTENNA__10330__S _11188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10851_ _19602_/Q _19440_/Q _18886_/Q _18656_/Q _10788_/S _10634_/A vssd1 vssd1 vccd1
+ vccd1 _10851_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17113__S _17119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _13570_/A _13570_/B _13584_/B _13570_/D vssd1 vssd1 vccd1 vccd1 _13571_/D
+ sky130_fd_sc_hd__nor4_1
X_10782_ _18432_/Q _09306_/A _09427_/A _10781_/X vssd1 vssd1 vccd1 vccd1 _12468_/A
+ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__17905__A1 _19754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12765__B _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _12791_/A _12751_/B _12791_/B vssd1 vssd1 vccd1 vccd1 _12602_/A sky130_fd_sc_hd__nor3_4
XANTENNA__11650__A0 _11070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _15240_/A vssd1 vssd1 vccd1 vccd1 _18682_/D sky130_fd_sc_hd__clkbuf_1
X_12452_ _12450_/Y _12451_/Y _12452_/S vssd1 vssd1 vccd1 vccd1 _12452_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15568__S _15568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ _18553_/Q _18552_/Q _18551_/Q _18550_/Q vssd1 vssd1 vccd1 vccd1 _11423_/A
+ sky130_fd_sc_hd__or4bb_2
X_15171_ _16673_/A vssd1 vssd1 vccd1 vccd1 _15171_/X sky130_fd_sc_hd__clkbuf_2
X_12383_ _12383_/A _14300_/B vssd1 vssd1 vccd1 vccd1 _12384_/B sky130_fd_sc_hd__nor2_1
XFILLER_126_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14122_ _13817_/X _14121_/X _14122_/S vssd1 vssd1 vccd1 vccd1 _14122_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11334_ _11372_/B _11584_/B _11585_/D _11333_/X vssd1 vssd1 vccd1 vccd1 _13521_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14053_ _14053_/A vssd1 vssd1 vccd1 vccd1 _18435_/D sky130_fd_sc_hd__clkbuf_1
X_18930_ _19642_/CLK _18930_/D vssd1 vssd1 vccd1 vccd1 _18930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11265_ _11242_/Y _11243_/X _11261_/X _11263_/Y _11264_/Y vssd1 vssd1 vccd1 vccd1
+ _11266_/D sky130_fd_sc_hd__a2111o_1
X_13004_ _13034_/A _13004_/B _13004_/C vssd1 vssd1 vccd1 vccd1 _18314_/D sky130_fd_sc_hd__nor3_1
X_10216_ _10210_/A _10213_/X _10215_/X _09988_/A vssd1 vssd1 vccd1 vccd1 _10216_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18861_ _19640_/CLK _18861_/D vssd1 vssd1 vccd1 vccd1 _18861_/Q sky130_fd_sc_hd__dfxtp_1
X_11196_ _09403_/A _11183_/X _11195_/X vssd1 vssd1 vccd1 vccd1 _11196_/X sky130_fd_sc_hd__a21o_2
XFILLER_95_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17812_ _15178_/X _19708_/Q _17816_/S vssd1 vssd1 vccd1 vccd1 _17813_/A sky130_fd_sc_hd__mux2_1
X_10147_ _10140_/Y _10142_/Y _10144_/Y _10146_/Y _09404_/A vssd1 vssd1 vccd1 vccd1
+ _10147_/X sky130_fd_sc_hd__o221a_1
XANTENNA__13458__A1 _13212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18792_ _19540_/CLK _18792_/D vssd1 vssd1 vccd1 vccd1 _18792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17743_ _18483_/Q _17743_/B vssd1 vssd1 vccd1 vccd1 _17743_/Y sky130_fd_sc_hd__nand2_1
X_14955_ _18478_/Q _18479_/Q _14955_/C vssd1 vssd1 vccd1 vccd1 _14979_/C sky130_fd_sc_hd__and3_1
X_10078_ _09783_/A _10075_/X _10077_/X vssd1 vssd1 vccd1 vccd1 _10078_/X sky130_fd_sc_hd__a21o_1
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_0_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13906_ _13753_/X _13667_/X _14278_/A _13905_/X vssd1 vssd1 vccd1 vccd1 _13906_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10240__S _10401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17674_ _18471_/Q _17674_/B vssd1 vssd1 vccd1 vccd1 _17675_/B sky130_fd_sc_hd__nand2_1
X_14886_ _14883_/Y _14884_/X _14885_/X _14838_/A _14999_/A vssd1 vssd1 vccd1 vccd1
+ _14887_/B sky130_fd_sc_hd__a221o_1
XANTENNA__12681__A2 _12665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19413_ _19706_/CLK _19413_/D vssd1 vssd1 vccd1 vccd1 _19413_/Q sky130_fd_sc_hd__dfxtp_1
X_16625_ _19268_/Q vssd1 vssd1 vccd1 vccd1 _16626_/A sky130_fd_sc_hd__clkbuf_1
X_13837_ _13745_/X _13964_/A _13836_/Y _13750_/X vssd1 vssd1 vccd1 vccd1 _13837_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__15080__A0 _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10119__S1 _09147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12969__B1 _12922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17023__S _17025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16556_ _19234_/Q _15564_/X _16558_/S vssd1 vssd1 vccd1 vccd1 _16557_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19344_ _19634_/CLK _19344_/D vssd1 vssd1 vccd1 vccd1 _19344_/Q sky130_fd_sc_hd__dfxtp_1
X_13768_ _13624_/X _13616_/X _13768_/S vssd1 vssd1 vccd1 vccd1 _13768_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09330__A _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12719_ _18279_/Q _12585_/A _12546_/A _13265_/A _12640_/A vssd1 vssd1 vccd1 vccd1
+ _12719_/X sky130_fd_sc_hd__a221o_1
X_15507_ _15590_/S vssd1 vssd1 vccd1 vccd1 _15520_/S sky130_fd_sc_hd__buf_2
X_16487_ _16487_/A vssd1 vssd1 vccd1 vccd1 _19203_/D sky130_fd_sc_hd__clkbuf_1
X_19275_ _19436_/CLK _19275_/D vssd1 vssd1 vccd1 vccd1 _19275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13699_ _13785_/A _13922_/B vssd1 vssd1 vccd1 vccd1 _13711_/B sky130_fd_sc_hd__nor2_4
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18226_ _18250_/A _18231_/C vssd1 vssd1 vccd1 vccd1 _18226_/Y sky130_fd_sc_hd__nor2_1
X_15438_ _15438_/A vssd1 vssd1 vccd1 vccd1 _18762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10195__B _12487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18157_ _18165_/A _18157_/B _18158_/B vssd1 vssd1 vccd1 vccd1 _19839_/D sky130_fd_sc_hd__nor3_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15369_ _18733_/Q _15178_/X _15373_/S vssd1 vssd1 vccd1 vccd1 _15370_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16163__A _16209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12691__A _13536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17108_ _16806_/X _19454_/Q _17108_/S vssd1 vssd1 vccd1 vccd1 _17109_/A sky130_fd_sc_hd__mux2_1
X_18088_ _18120_/A _18088_/B _18088_/C vssd1 vssd1 vccd1 vccd1 _19815_/D sky130_fd_sc_hd__nor3_1
X_09930_ _18609_/Q _19298_/Q _09955_/A vssd1 vssd1 vccd1 vccd1 _09930_/X sky130_fd_sc_hd__mux2_1
X_17039_ _19423_/Q _16705_/X _17047_/S vssd1 vssd1 vccd1 vccd1 _17040_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09861_ _09861_/A _09861_/B vssd1 vssd1 vccd1 vccd1 _09861_/X sky130_fd_sc_hd__or2_1
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15507__A _15590_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09792_ _10074_/A vssd1 vssd1 vccd1 vccd1 _09992_/A sky130_fd_sc_hd__clkbuf_2
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09748__S0 _09734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12672__A2 _13235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15071__A0 _18457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13621__A1 _12180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09240__A _09856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09920__S0 _09914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10386__A _10400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09226_ _09459_/A vssd1 vssd1 vccd1 vccd1 _09227_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14177__A2 _14176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13697__A _13720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09157_ _09643_/S vssd1 vssd1 vccd1 vccd1 _11157_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_148_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15126__B2 _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09088_ _09088_/A vssd1 vssd1 vccd1 vccd1 _11339_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13137__B1 _14673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14885__A0 _18441_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13688__A1 _14093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12104__A1_N _14555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11050_ _18586_/Q _19275_/Q _11050_/S vssd1 vssd1 vccd1 vccd1 _11050_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10001_ _09992_/X _09994_/X _09998_/X _10000_/X _09249_/X vssd1 vssd1 vccd1 vccd1
+ _10001_/X sky130_fd_sc_hd__a221o_2
XFILLER_131_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17823__A0 _15194_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17108__S _17108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15417__A _15485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16012__S _16016_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09415__A _09892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16947__S _16953_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11156__S _11156_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14740_ _16752_/A vssd1 vssd1 vccd1 vccd1 _14740_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11952_ _11952_/A vssd1 vssd1 vccd1 vccd1 _11954_/A sky130_fd_sc_hd__inv_2
XFILLER_123_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10903_ _18428_/Q vssd1 vssd1 vccd1 vccd1 _10903_/Y sky130_fd_sc_hd__inv_2
X_14671_ input49/X _14640_/X _14643_/X _14570_/A vssd1 vssd1 vccd1 vccd1 _15958_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11883_ _11880_/A _11882_/Y _12165_/S vssd1 vssd1 vccd1 vccd1 _11883_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16410_ _16410_/A vssd1 vssd1 vccd1 vccd1 _19169_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11680__A _16212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13622_ _13622_/A vssd1 vssd1 vccd1 vccd1 _14057_/B sky130_fd_sc_hd__buf_2
X_17390_ _17390_/A vssd1 vssd1 vccd1 vccd1 _19564_/D sky130_fd_sc_hd__clkbuf_1
X_10834_ _09273_/A _10823_/X _10833_/X _09280_/A _18430_/Q vssd1 vssd1 vccd1 vccd1
+ _10834_/X sky130_fd_sc_hd__a32o_2
XANTENNA__09816__B1 _09320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12495__B _12495_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16341_ _16341_/A vssd1 vssd1 vccd1 vccd1 _19139_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10426__A1 _09689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13553_ _09109_/Y _13536_/X _13537_/X _14802_/B vssd1 vssd1 vccd1 vccd1 _13554_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_160_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10765_ _19635_/Q _19052_/Q _19089_/Q _18695_/Q _10650_/S _09482_/A vssd1 vssd1 vccd1
+ vccd1 _10765_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10296__A _18442_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19060_ _19579_/CLK _19060_/D vssd1 vssd1 vccd1 vccd1 _19060_/Q sky130_fd_sc_hd__dfxtp_1
X_12504_ _12504_/A _12505_/B vssd1 vssd1 vccd1 vccd1 _12504_/Y sky130_fd_sc_hd__nor2_1
X_16272_ _16272_/A vssd1 vssd1 vccd1 vccd1 _19108_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_190_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19608_/CLK sky130_fd_sc_hd__clkbuf_16
X_13484_ _18401_/Q _12617_/B _13486_/S vssd1 vssd1 vccd1 vccd1 _13485_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10696_ _11065_/A vssd1 vssd1 vccd1 vccd1 _10791_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18011_ _19789_/Q _19788_/Q _18011_/C vssd1 vssd1 vccd1 vccd1 _18014_/B sky130_fd_sc_hd__and3_1
X_15223_ _16725_/A vssd1 vssd1 vccd1 vccd1 _15223_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15298__S _15300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12435_ _12219_/S _12433_/X _12451_/B _11847_/X vssd1 vssd1 vccd1 vccd1 _12435_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_139_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15154_ _15154_/A vssd1 vssd1 vccd1 vccd1 _18655_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_0_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12366_ _18377_/Q vssd1 vssd1 vccd1 vccd1 _13388_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15117__B2 _11139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_153_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14105_ _14122_/S _13854_/X _14104_/X vssd1 vssd1 vccd1 vccd1 _14105_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_4_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11317_ _11317_/A vssd1 vssd1 vccd1 vccd1 _11365_/A sky130_fd_sc_hd__inv_2
XFILLER_126_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14930__S _14941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17807__A _17853_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15085_ _15085_/A vssd1 vssd1 vccd1 vccd1 _18620_/D sky130_fd_sc_hd__clkbuf_1
X_12297_ _18374_/Q vssd1 vssd1 vccd1 vccd1 _13352_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13679__A1 _14074_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14036_ _13972_/Y _14035_/Y _14036_/S vssd1 vssd1 vccd1 vccd1 _14036_/X sky130_fd_sc_hd__mux2_1
X_18913_ _18982_/CLK _18913_/D vssd1 vssd1 vccd1 vccd1 _18913_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output75_A _11956_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11248_ _11248_/A _11248_/B _11248_/C vssd1 vssd1 vccd1 vccd1 _11248_/Y sky130_fd_sc_hd__nand3_1
XFILLER_68_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17814__A0 _15181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12351__A1 _18517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18844_ _19643_/CLK _18844_/D vssd1 vssd1 vccd1 vccd1 _18844_/Q sky130_fd_sc_hd__dfxtp_1
X_11179_ _19529_/Q _19143_/Q _19593_/Q _18749_/Q _09729_/S _09728_/A vssd1 vssd1 vccd1
+ vccd1 _11180_/B sky130_fd_sc_hd__mux4_1
XFILLER_110_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18775_ _19555_/CLK _18775_/D vssd1 vssd1 vccd1 vccd1 _18775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12103__A1 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15987_ _15987_/A vssd1 vssd1 vccd1 vccd1 _18992_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15761__S _15769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17726_ _19680_/Q _17708_/X _17722_/Y _17725_/X vssd1 vssd1 vccd1 vccd1 _19680_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_48_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14938_ _14934_/X _14936_/Y _14937_/Y vssd1 vssd1 vccd1 vccd1 _16702_/A sky130_fd_sc_hd__a21oi_4
XFILLER_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10665__A1 _10366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_143_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _18982_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17657_ _17667_/C _17657_/B vssd1 vssd1 vccd1 vccd1 _17657_/Y sky130_fd_sc_hd__nand2_2
X_14869_ _14869_/A vssd1 vssd1 vccd1 vccd1 _18599_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11590__A _11618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16608_ _16608_/A vssd1 vssd1 vccd1 vccd1 _19259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_78_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17588_ _19652_/Q _16819_/A _17590_/S vssd1 vssd1 vccd1 vccd1 _17589_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19327_ _19553_/CLK _19327_/D vssd1 vssd1 vccd1 vccd1 _19327_/Q sky130_fd_sc_hd__dfxtp_1
X_16539_ _19226_/Q _15538_/X _16547_/S vssd1 vssd1 vccd1 vccd1 _16540_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_158_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _18853_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11090__A1 _09695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15356__A1 _15159_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19258_ _19580_/CLK _19258_/D vssd1 vssd1 vccd1 vccd1 _19258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18209_ _19857_/Q _18214_/B _12948_/X vssd1 vssd1 vccd1 vccd1 _18210_/B sky130_fd_sc_hd__o21ai_1
XFILLER_148_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19189_ _19706_/CLK _19189_/D vssd1 vssd1 vccd1 vccd1 _19189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15108__A1 _18632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15108__B2 _11130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09913_ _19330_/Q vssd1 vssd1 vccd1 vccd1 _09913_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12342__A1 _12193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17805__A0 _15168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09844_ _18874_/Q _19332_/Q _09911_/S vssd1 vssd1 vccd1 vccd1 _09844_/X sky130_fd_sc_hd__mux2_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09235__A _09856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09775_ _09770_/X _09771_/X _09908_/A vssd1 vssd1 vccd1 vccd1 _09775_/X sky130_fd_sc_hd__a21o_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16068__A _16135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10751__S1 _10670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15595__A1 _15487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10550_ _10622_/A _10550_/B vssd1 vssd1 vccd1 vccd1 _10550_/X sky130_fd_sc_hd__or2_1
XFILLER_168_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09209_ _09209_/A vssd1 vssd1 vccd1 vccd1 _09210_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_154_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10481_ _11099_/A _10478_/X _10480_/X _09227_/A vssd1 vssd1 vccd1 vccd1 _10481_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12476__A_N _12472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12220_ _12214_/Y _12219_/X _13529_/B vssd1 vssd1 vccd1 vccd1 _12220_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10267__S0 _11156_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11659__B _11788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15846__S _15852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12151_ _13316_/A _12169_/C _12150_/Y vssd1 vssd1 vccd1 vccd1 _12151_/X sky130_fd_sc_hd__o21a_1
XFILLER_151_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10019__S0 _09782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11102_ _11102_/A _11102_/B vssd1 vssd1 vccd1 vccd1 _11102_/X sky130_fd_sc_hd__or2_1
XFILLER_151_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12082_ _14155_/A _12082_/B vssd1 vssd1 vccd1 vccd1 _12085_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13530__B1 _14519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15910_ _15910_/A vssd1 vssd1 vccd1 vccd1 _18957_/D sky130_fd_sc_hd__clkbuf_1
X_11033_ _10956_/A _11032_/X _09223_/A vssd1 vssd1 vccd1 vccd1 _11033_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16890_ _16890_/A vssd1 vssd1 vccd1 vccd1 _19357_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09145__A _09145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15841_ _14879_/X _18927_/Q _15841_/S vssd1 vssd1 vccd1 vccd1 _15842_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14986__A _16819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_60_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19718_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__15581__S _15584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18560_ _18585_/CLK _18560_/D vssd1 vssd1 vccd1 vccd1 _18560_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _18308_/Q _18307_/Q _18309_/Q _12984_/D vssd1 vssd1 vccd1 vccd1 _12995_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_18_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15772_ _14889_/X _18896_/Q _15780_/S vssd1 vssd1 vccd1 vccd1 _15773_/A sky130_fd_sc_hd__mux2_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ _17511_/A vssd1 vssd1 vccd1 vccd1 _19617_/D sky130_fd_sc_hd__clkbuf_1
X_11935_ _11930_/Y _11933_/X _11934_/X _11560_/X vssd1 vssd1 vccd1 vccd1 _11935_/X
+ sky130_fd_sc_hd__o211a_1
X_14723_ _14714_/X _18586_/Q _14762_/S vssd1 vssd1 vccd1 vccd1 _14724_/A sky130_fd_sc_hd__mux2_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18491_ _18623_/CLK _18491_/D vssd1 vssd1 vccd1 vccd1 _18491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10742__S1 _10670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17442_ _16816_/X _19587_/Q _17446_/S vssd1 vssd1 vccd1 vccd1 _17443_/A sky130_fd_sc_hd__mux2_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ _14654_/A _17777_/B vssd1 vssd1 vccd1 vccd1 _14655_/A sky130_fd_sc_hd__and2_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _11970_/A _11866_/B vssd1 vssd1 vccd1 vccd1 _11867_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_75_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19806_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13597__A0 _14111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13605_ _13643_/A vssd1 vssd1 vccd1 vccd1 _13685_/S sky130_fd_sc_hd__buf_2
X_10817_ _10813_/X _10815_/X _10816_/X _11041_/A _09208_/A vssd1 vssd1 vccd1 vccd1
+ _10823_/B sky130_fd_sc_hd__o221a_1
X_17373_ _17373_/A vssd1 vssd1 vccd1 vccd1 _19556_/D sky130_fd_sc_hd__clkbuf_1
X_14585_ _14585_/A vssd1 vssd1 vccd1 vccd1 _14585_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_159_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11797_ _11768_/A _11766_/X _11767_/A vssd1 vssd1 vccd1 vccd1 _11823_/B sky130_fd_sc_hd__a21o_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16706__A _16722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19112_ _19724_/CLK _19112_/D vssd1 vssd1 vccd1 vccd1 _19112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16324_ _16324_/A vssd1 vssd1 vccd1 vccd1 _19131_/D sky130_fd_sc_hd__clkbuf_1
X_13536_ _13536_/A vssd1 vssd1 vccd1 vccd1 _13536_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10748_ _09209_/A _10743_/X _10745_/X _10747_/X _10568_/A vssd1 vssd1 vccd1 vccd1
+ _10748_/X sky130_fd_sc_hd__a221o_2
XANTENNA__11072__B2 _12463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16255_ _16093_/X _19101_/Q _16257_/S vssd1 vssd1 vccd1 vccd1 _16256_/A sky130_fd_sc_hd__mux2_1
X_19043_ _19725_/CLK _19043_/D vssd1 vssd1 vccd1 vccd1 _19043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13467_ _18393_/Q _13259_/X _13475_/S vssd1 vssd1 vccd1 vccd1 _13468_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10679_ _19410_/Q _19186_/Q _19703_/Q _19154_/Q _10860_/S _09139_/A vssd1 vssd1 vccd1
+ vccd1 _10679_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13130__A _13130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15206_ _15206_/A vssd1 vssd1 vccd1 vccd1 _18671_/D sky130_fd_sc_hd__clkbuf_1
X_12418_ _14587_/A _13525_/A _12345_/X _12504_/A vssd1 vssd1 vccd1 vccd1 _12419_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_16186_ _16099_/X _19066_/Q _16194_/S vssd1 vssd1 vccd1 vccd1 _16187_/A sky130_fd_sc_hd__mux2_1
X_13398_ _18647_/Q _13398_/B vssd1 vssd1 vccd1 vccd1 _13398_/X sky130_fd_sc_hd__or2_1
XFILLER_154_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15137_ _16503_/A vssd1 vssd1 vccd1 vccd1 _16847_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_99_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17537__A _17605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12349_ _13712_/A _14274_/B _12327_/B vssd1 vssd1 vccd1 vccd1 _12350_/B sky130_fd_sc_hd__a21o_1
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19549_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_141_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15068_ _15068_/A vssd1 vssd1 vccd1 vccd1 _18616_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14019_ _14001_/Y _14018_/Y _14019_/S vssd1 vssd1 vccd1 vccd1 _14019_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12324__B2 _12500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10335__B1 _09394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18827_ _19543_/CLK _18827_/D vssd1 vssd1 vccd1 vccd1 _18827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_28_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19165_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09560_ _18782_/Q _19011_/Q _18942_/Q _19240_/Q _09700_/A _09642_/A vssd1 vssd1 vccd1
+ vccd1 _09561_/B sky130_fd_sc_hd__mux4_1
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18758_ _19569_/CLK _18758_/D vssd1 vssd1 vccd1 vccd1 _18758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12627__A2 _13236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11835__A0 _11834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17709_ _18477_/Q _17710_/B vssd1 vssd1 vccd1 vccd1 _17720_/C sky130_fd_sc_hd__or2_1
X_09491_ _10500_/A vssd1 vssd1 vccd1 vccd1 _10511_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18689_ _19632_/CLK _18689_/D vssd1 vssd1 vccd1 vccd1 _18689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13305__A _18634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10497__S0 _10450_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15501__A1 _15500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11495__A _11511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09827_ _10140_/A vssd1 vssd1 vccd1 vccd1 _10042_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14068__A1 _11926_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16497__S _16497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10972__S1 _10920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09758_ _10094_/A vssd1 vssd1 vccd1 vccd1 _10076_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_58_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_101_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _09689_/A vssd1 vssd1 vccd1 vccd1 _09689_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13291__A2 _12735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _11720_/A _11720_/B vssd1 vssd1 vccd1 vccd1 _11820_/B sky130_fd_sc_hd__nor2_2
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _11652_/A _13665_/A vssd1 vssd1 vccd1 vccd1 _11653_/A sky130_fd_sc_hd__and2_1
XFILLER_14_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10602_ _19251_/Q _19022_/Q _18953_/Q _19347_/Q _10605_/S _10366_/A vssd1 vssd1 vccd1
+ vccd1 _10603_/B sky130_fd_sc_hd__mux4_1
XFILLER_11_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10488__S0 _10389_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14370_ _18468_/Q _18500_/Q _14381_/S vssd1 vssd1 vccd1 vccd1 _14371_/A sky130_fd_sc_hd__mux2_1
X_11582_ _18561_/Q _11556_/A _11576_/X _11581_/Y vssd1 vssd1 vccd1 vccd1 _11688_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_13321_ _13365_/A vssd1 vssd1 vccd1 vccd1 _13352_/B sky130_fd_sc_hd__clkbuf_2
X_10533_ _19607_/Q _19445_/Q _18891_/Q _18661_/Q _10558_/S _10367_/A vssd1 vssd1 vccd1
+ vccd1 _10534_/B sky130_fd_sc_hd__mux4_1
XFILLER_7_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16960__S _16964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16040_ _16039_/X _19015_/Q _16049_/S vssd1 vssd1 vccd1 vccd1 _16041_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12003__B1 _17878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13252_ _19669_/Q _13251_/X _12768_/X _18393_/Q vssd1 vssd1 vccd1 vccd1 _13253_/B
+ sky130_fd_sc_hd__a22o_1
X_10464_ _10477_/A _10464_/B vssd1 vssd1 vccd1 vccd1 _10464_/X sky130_fd_sc_hd__or2_1
XFILLER_170_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12203_ _12491_/C _12226_/A _12202_/X vssd1 vssd1 vccd1 vccd1 _14216_/A sky130_fd_sc_hd__o21ai_4
XFILLER_142_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13183_ _18354_/Q _13183_/B vssd1 vssd1 vccd1 vccd1 _13183_/X sky130_fd_sc_hd__or2_1
XFILLER_135_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10395_ _10395_/A vssd1 vssd1 vccd1 vccd1 _10438_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12134_ _12177_/A vssd1 vssd1 vccd1 vccd1 _12328_/A sky130_fd_sc_hd__buf_2
XFILLER_89_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17991_ _17991_/A _17997_/C vssd1 vssd1 vccd1 vccd1 _17991_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19730_ _19732_/CLK _19730_/D vssd1 vssd1 vccd1 vccd1 _19730_/Q sky130_fd_sc_hd__dfxtp_2
X_16942_ _16774_/X _19380_/Q _16942_/S vssd1 vssd1 vccd1 vccd1 _16943_/A sky130_fd_sc_hd__mux2_1
X_12065_ _12040_/A _12040_/B _12036_/A vssd1 vssd1 vccd1 vccd1 _12066_/B sky130_fd_sc_hd__a21oi_2
XFILLER_145_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11016_ _11062_/A _11016_/B vssd1 vssd1 vccd1 vccd1 _11016_/X sky130_fd_sc_hd__or2_1
X_19661_ _19689_/CLK _19661_/D vssd1 vssd1 vccd1 vccd1 _19661_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__13109__B _13536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16873_ _16873_/A vssd1 vssd1 vccd1 vccd1 _19349_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10332__A3 _19354_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18612_ _19591_/CLK _18612_/D vssd1 vssd1 vccd1 vccd1 _18612_/Q sky130_fd_sc_hd__dfxtp_1
X_15824_ _14782_/X _18919_/Q _15830_/S vssd1 vssd1 vccd1 vccd1 _15825_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15605__A _15662_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19592_ _19592_/CLK _19592_/D vssd1 vssd1 vccd1 vccd1 _19592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18543_ _19732_/CLK _18543_/D vssd1 vssd1 vccd1 vccd1 _18543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ _12972_/A _14638_/A vssd1 vssd1 vccd1 vccd1 _18303_/D sky130_fd_sc_hd__nor2_1
X_15755_ _15755_/A vssd1 vssd1 vccd1 vccd1 _18888_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10715__S1 _09352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16756__A0 _16755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11918_ _11918_/A _13622_/A vssd1 vssd1 vccd1 vccd1 _11919_/B sky130_fd_sc_hd__or2_1
X_14706_ _19079_/Q vssd1 vssd1 vccd1 vccd1 _14825_/A sky130_fd_sc_hd__inv_2
XFILLER_61_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18474_ _19079_/CLK _18474_/D vssd1 vssd1 vccd1 vccd1 _18474_/Q sky130_fd_sc_hd__dfxtp_1
X_12898_ _18278_/Q _12894_/C _12897_/Y vssd1 vssd1 vccd1 vccd1 _18278_/D sky130_fd_sc_hd__o21a_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15686_ _18858_/Q _15519_/X _15686_/S vssd1 vssd1 vccd1 vccd1 _15687_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _17425_/A vssd1 vssd1 vccd1 vccd1 _19579_/D sky130_fd_sc_hd__clkbuf_1
X_11849_ _11849_/A _19735_/Q _12095_/B vssd1 vssd1 vccd1 vccd1 _11850_/A sky130_fd_sc_hd__and3_1
X_14637_ input37/X _14593_/X _14597_/X _14543_/A vssd1 vssd1 vccd1 vccd1 _14638_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ _14568_/A _14580_/B vssd1 vssd1 vccd1 vccd1 _14568_/X sky130_fd_sc_hd__or2_1
XANTENNA__10479__S0 _09449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17356_ _17356_/A vssd1 vssd1 vccd1 vccd1 _19548_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12683__B _12683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16307_ _16064_/X _19124_/Q _16307_/S vssd1 vssd1 vccd1 vccd1 _16308_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17181__A0 _18438_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13519_ _11313_/D _11552_/B _11551_/Y _09113_/B vssd1 vssd1 vccd1 vccd1 _13520_/C
+ sky130_fd_sc_hd__o2bb2a_1
X_14499_ _14499_/A vssd1 vssd1 vccd1 vccd1 _18519_/D sky130_fd_sc_hd__clkbuf_1
X_17287_ _19518_/Q _16696_/X _17291_/S vssd1 vssd1 vccd1 vccd1 _17288_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19026_ _19710_/CLK _19026_/D vssd1 vssd1 vccd1 vccd1 _19026_/Q sky130_fd_sc_hd__dfxtp_1
X_16238_ _16067_/X _19093_/Q _16246_/S vssd1 vssd1 vccd1 vccd1 _16239_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16169_ _16169_/A vssd1 vssd1 vccd1 vccd1 _19058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10859__A1 _09629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19859_ _19859_/CLK _19859_/D vssd1 vssd1 vccd1 vccd1 _19859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10323__A3 _10322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09612_ _10177_/A _09612_/B vssd1 vssd1 vccd1 vccd1 _09612_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16110__S _16113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_15_0_clock_A clkbuf_3_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09513__A _10887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09543_ _09643_/S vssd1 vssd1 vccd1 vccd1 _09793_/A sky130_fd_sc_hd__buf_4
XFILLER_52_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14470__A1 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17730__A _17730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09474_ _10764_/A vssd1 vssd1 vccd1 vccd1 _10591_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16747__A0 _16743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12874__A _12904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14222__A1 _18447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14222__B2 _14221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10244__C1 _10400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10890__S0 _11050_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10180_ _09414_/A _10173_/Y _10175_/Y _10177_/Y _10179_/Y vssd1 vssd1 vccd1 vccd1
+ _10180_/X sky130_fd_sc_hd__o32a_1
XFILLER_78_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10945__S1 _09481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13870_ _13870_/A _13870_/B vssd1 vssd1 vccd1 vccd1 _14115_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12821_ _18256_/Q _12821_/B _12821_/C vssd1 vssd1 vccd1 vccd1 _12822_/C sky130_fd_sc_hd__and3_1
XFILLER_62_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14461__A1 _17878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ _12752_/A vssd1 vssd1 vccd1 vccd1 _12753_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15540_ _18800_/Q _15538_/X _15552_/S vssd1 vssd1 vccd1 vccd1 _15541_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _11702_/B _11703_/B vssd1 vssd1 vccd1 vccd1 _11704_/B sky130_fd_sc_hd__and2b_1
XFILLER_42_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15471_ _15471_/A vssd1 vssd1 vccd1 vccd1 _18777_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12712_/A _12683_/B vssd1 vssd1 vccd1 vccd1 _12683_/Y sky130_fd_sc_hd__nor2_2
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _19489_/Q _17208_/X _17223_/S vssd1 vssd1 vccd1 vccd1 _17211_/A sky130_fd_sc_hd__mux2_1
X_14422_ _14422_/A vssd1 vssd1 vccd1 vccd1 _18486_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11634_ _11835_/S vssd1 vssd1 vccd1 vccd1 _12173_/A sky130_fd_sc_hd__buf_2
X_18190_ _19850_/Q _18191_/C _19851_/Q vssd1 vssd1 vccd1 vccd1 _18192_/B sky130_fd_sc_hd__a21oi_1
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11122__S1 _10451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17141_ _19469_/Q _17136_/X _17155_/S vssd1 vssd1 vccd1 vccd1 _17142_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17786__S _17794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14353_ _14353_/A vssd1 vssd1 vccd1 vccd1 _18462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11565_ _11565_/A _11565_/B _11565_/C vssd1 vssd1 vccd1 vccd1 _11749_/A sky130_fd_sc_hd__and3_2
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13304_ _19775_/Q _13123_/A _13300_/X _13303_/X vssd1 vssd1 vccd1 vccd1 _13305_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_10_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17072_ _17072_/A vssd1 vssd1 vccd1 vccd1 _19437_/D sky130_fd_sc_hd__clkbuf_1
X_10516_ _10640_/A _10516_/B vssd1 vssd1 vccd1 vccd1 _10516_/X sky130_fd_sc_hd__or2_1
XFILLER_171_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14284_ _14284_/A _14319_/B vssd1 vssd1 vccd1 vccd1 _14284_/Y sky130_fd_sc_hd__nor2_1
X_11496_ _11664_/B _11519_/C _11664_/C vssd1 vssd1 vccd1 vccd1 _11506_/A sky130_fd_sc_hd__or3_1
XFILLER_171_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13235_ _13235_/A vssd1 vssd1 vccd1 vccd1 _13235_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16023_ _15033_/X _19009_/Q _16027_/S vssd1 vssd1 vccd1 vccd1 _16024_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10447_ _10447_/A _10447_/B vssd1 vssd1 vccd1 vccd1 _10447_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14504__A _18225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10002__A2 _09990_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17466__A1 _16639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ _13166_/A _13183_/B vssd1 vssd1 vccd1 vccd1 _13166_/X sky130_fd_sc_hd__or2_1
X_10378_ _18831_/Q _19385_/Q _19547_/Q _18799_/Q _09448_/S _10349_/A vssd1 vssd1 vccd1
+ vccd1 _10379_/B sky130_fd_sc_hd__mux4_1
XFILLER_151_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12117_ _19744_/Q _12117_/B _12117_/C vssd1 vssd1 vccd1 vccd1 _12144_/C sky130_fd_sc_hd__and3_1
XANTENNA__10553__A3 _10552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17974_ _17991_/A _17979_/C vssd1 vssd1 vccd1 vccd1 _17974_/Y sky130_fd_sc_hd__nor2_1
X_13097_ _17781_/A vssd1 vssd1 vccd1 vccd1 _14612_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_112_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17218__A1 _12757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19713_ _19713_/CLK _19713_/D vssd1 vssd1 vccd1 vccd1 _19713_/Q sky130_fd_sc_hd__dfxtp_1
X_12048_ _12098_/B _12045_/X _12047_/Y vssd1 vssd1 vccd1 vccd1 _12048_/Y sky130_fd_sc_hd__a21oi_1
X_16925_ _16749_/X _19372_/Q _16931_/S vssd1 vssd1 vccd1 vccd1 _16926_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10936__S1 _09352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19644_ _19714_/CLK _19644_/D vssd1 vssd1 vccd1 vccd1 _19644_/Q sky130_fd_sc_hd__dfxtp_1
X_16856_ _19342_/Q _16651_/X _16858_/S vssd1 vssd1 vccd1 vccd1 _16857_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09333__A _09969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15807_ _15807_/A vssd1 vssd1 vccd1 vccd1 _18912_/D sky130_fd_sc_hd__clkbuf_1
X_19575_ _19639_/CLK _19575_/D vssd1 vssd1 vccd1 vccd1 _19575_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16865__S _16869_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16787_ _16787_/A vssd1 vssd1 vccd1 vccd1 _16787_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14452__A1 _11901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13999_ _13995_/X _13998_/Y _13999_/S vssd1 vssd1 vccd1 vccd1 _13999_/X sky130_fd_sc_hd__mux2_2
XFILLER_46_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18526_ _18567_/CLK _18526_/D vssd1 vssd1 vccd1 vccd1 _18526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15738_ _15806_/S vssd1 vssd1 vccd1 vccd1 _15747_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_80_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18457_ _19695_/CLK _18457_/D vssd1 vssd1 vccd1 vccd1 _18457_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12694__A _13042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15669_ _18850_/Q _15494_/X _15675_/S vssd1 vssd1 vccd1 vccd1 _15670_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17408_ _17408_/A vssd1 vssd1 vccd1 vccd1 _19571_/D sky130_fd_sc_hd__clkbuf_1
X_09190_ _09190_/A vssd1 vssd1 vccd1 vccd1 _09190_/X sky130_fd_sc_hd__buf_2
X_18388_ _19791_/CLK _18388_/D vssd1 vssd1 vccd1 vccd1 _18388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17154__A0 _10810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17339_ _16771_/X _19541_/Q _17341_/S vssd1 vssd1 vccd1 vccd1 _17340_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10418__S _10465_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10872__S0 _10664_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19009_ _19579_/CLK _19009_/D vssd1 vssd1 vccd1 vccd1 _19009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15944__S _15946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10153__S _10153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12869__A _18173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11492__B _14587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14443__A1 _19732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09526_ _19531_/Q _19145_/Q _19595_/Q _18751_/Q _10242_/S _09501_/A vssd1 vssd1 vccd1
+ vccd1 _09527_/B sky130_fd_sc_hd__mux4_1
XFILLER_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09457_ _18783_/Q _19012_/Q _18943_/Q _19241_/Q _10540_/S _09141_/A vssd1 vssd1 vccd1
+ vccd1 _09458_/B sky130_fd_sc_hd__mux4_1
XFILLER_52_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09897__B _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09388_ _09421_/A _09372_/X _09387_/X vssd1 vssd1 vccd1 vccd1 _09388_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10217__C1 _09248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10328__S _10328_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ _18580_/Q _18579_/Q _18568_/Q _18567_/Q vssd1 vssd1 vccd1 vccd1 _11356_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_153_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ _19516_/Q _19130_/Q _19580_/Q _18736_/Q _09701_/S _09555_/X vssd1 vssd1 vccd1
+ vccd1 _10302_/B sky130_fd_sc_hd__mux4_1
X_11281_ _11501_/B _11285_/B vssd1 vssd1 vccd1 vccd1 _11281_/Y sky130_fd_sc_hd__nand2_1
XFILLER_106_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14324__A _14324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13020_ _18318_/Q _13016_/C _13019_/Y vssd1 vssd1 vccd1 vccd1 _18318_/D sky130_fd_sc_hd__o21a_1
XFILLER_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13182__B2 _18623_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10232_ _19646_/Q _19063_/Q _19100_/Q _18706_/Q _10230_/X _11111_/A vssd1 vssd1 vccd1
+ vccd1 _10232_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11667__B _11667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11193__B1 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14043__B _14045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17635__A _17693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10163_ _10167_/A _10163_/B vssd1 vssd1 vccd1 vccd1 _10163_/X sky130_fd_sc_hd__or2_1
XFILLER_126_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input37_A io_ibus_inst[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ _10094_/A vssd1 vssd1 vccd1 vccd1 _10094_/X sky130_fd_sc_hd__buf_2
X_14971_ _14838_/X _14970_/X _14898_/X vssd1 vssd1 vccd1 vccd1 _14971_/Y sky130_fd_sc_hd__a21oi_2
X_16710_ _19296_/Q _16709_/X _16719_/S vssd1 vssd1 vccd1 vccd1 _16711_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11040__S0 _10959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13922_ _13922_/A _13922_/B vssd1 vssd1 vccd1 vccd1 _13942_/A sky130_fd_sc_hd__nor2_2
XFILLER_59_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09784__S1 _09783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17690_ _18474_/Q _17691_/B vssd1 vssd1 vccd1 vccd1 _17701_/C sky130_fd_sc_hd__or2_1
XFILLER_19_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09153__A _10605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16641_ _16722_/A vssd1 vssd1 vccd1 vccd1 _16741_/S sky130_fd_sc_hd__buf_8
XFILLER_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13853_ _13966_/S _13776_/X _13813_/Y vssd1 vssd1 vccd1 vccd1 _13853_/X sky130_fd_sc_hd__o21a_1
XFILLER_90_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10299__A _10299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12804_ _12808_/B _18250_/B _12803_/Y vssd1 vssd1 vccd1 vccd1 _18252_/D sky130_fd_sc_hd__o21a_1
X_19360_ _19717_/CLK _19360_/D vssd1 vssd1 vccd1 vccd1 _19360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16572_ _16572_/A vssd1 vssd1 vccd1 vccd1 _19241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09536__S1 _09144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13784_ _14097_/A vssd1 vssd1 vccd1 vccd1 _13784_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10996_ _10996_/A _10996_/B vssd1 vssd1 vccd1 vccd1 _10996_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18311_ _19798_/CLK _18311_/D vssd1 vssd1 vccd1 vccd1 _18311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15523_ _15590_/S vssd1 vssd1 vccd1 vccd1 _15536_/S sky130_fd_sc_hd__buf_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _12735_/A vssd1 vssd1 vccd1 vccd1 _12736_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19291_ _19612_/CLK _19291_/D vssd1 vssd1 vccd1 vccd1 _19291_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18242_ _18242_/A vssd1 vssd1 vccd1 vccd1 _18247_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12666_ _19763_/Q _12666_/B vssd1 vssd1 vccd1 vccd1 _12666_/X sky130_fd_sc_hd__or2_1
XFILLER_124_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _15454_/A vssd1 vssd1 vccd1 vccd1 _18769_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10208__C1 _09134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17136__A0 _11046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11617_ _13625_/A _11940_/A _13769_/S vssd1 vssd1 vccd1 vccd1 _11622_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__11307__B1_N input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14405_ _14405_/A vssd1 vssd1 vccd1 vccd1 _18480_/D sky130_fd_sc_hd__clkbuf_1
X_18173_ _18173_/A vssd1 vssd1 vccd1 vccd1 _18249_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12597_ _12577_/X _12579_/Y _12594_/X _12596_/X _18636_/Q vssd1 vssd1 vccd1 vccd1
+ _12598_/B sky130_fd_sc_hd__a32o_4
X_15385_ _15385_/A vssd1 vssd1 vccd1 vccd1 _18740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17124_ _16829_/X _19461_/Q _17130_/S vssd1 vssd1 vccd1 vccd1 _17125_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14336_ _13696_/X _14150_/A _14335_/X _13832_/A vssd1 vssd1 vccd1 vccd1 _14336_/X
+ sky130_fd_sc_hd__a211o_1
X_11548_ _15071_/S vssd1 vssd1 vccd1 vccd1 _15018_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_144_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14267_ _14182_/A _14264_/X _14266_/Y _13950_/A vssd1 vssd1 vccd1 vccd1 _14267_/X
+ sky130_fd_sc_hd__a31o_1
X_17055_ _17055_/A vssd1 vssd1 vccd1 vccd1 _19430_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11479_ _11479_/A vssd1 vssd1 vccd1 vccd1 _13521_/A sky130_fd_sc_hd__inv_2
XFILLER_100_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13218_ _13248_/A _18627_/Q vssd1 vssd1 vccd1 vccd1 _13218_/Y sky130_fd_sc_hd__nand2_1
X_16006_ _16006_/A vssd1 vssd1 vccd1 vccd1 _19001_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14198_ _18445_/Q _14120_/X _14197_/X vssd1 vssd1 vccd1 vccd1 _18445_/D sky130_fd_sc_hd__o21a_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13149_ _13121_/X _13140_/Y _13148_/X _13135_/X _18620_/Q vssd1 vssd1 vccd1 vccd1
+ _13149_/X sky130_fd_sc_hd__a32o_4
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _19770_/Q _19769_/Q _19768_/Q _17957_/D vssd1 vssd1 vccd1 vccd1 _17963_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_140_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11593__A _11593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16908_ _16908_/A vssd1 vssd1 vccd1 vccd1 _19365_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15065__A _16737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11031__S0 _10959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17888_ _17890_/A _17888_/B vssd1 vssd1 vccd1 vccd1 _17889_/A sky130_fd_sc_hd__and2_1
XFILLER_93_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19627_ _19726_/CLK _19627_/D vssd1 vssd1 vccd1 vccd1 _19627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16839_ _16838_/X _19336_/Q _16839_/S vssd1 vssd1 vccd1 vccd1 _16840_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19558_ _19590_/CLK _19558_/D vssd1 vssd1 vccd1 vccd1 _19558_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_148_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09311_ _10728_/A vssd1 vssd1 vccd1 vccd1 _10793_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18509_ _18509_/CLK _18509_/D vssd1 vssd1 vccd1 vccd1 _18509_/Q sky130_fd_sc_hd__dfxtp_1
X_19489_ _19496_/CLK _19489_/D vssd1 vssd1 vccd1 vccd1 _19489_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10998__B1 _09223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09242_ _19695_/Q vssd1 vssd1 vccd1 vccd1 _09243_/A sky130_fd_sc_hd__inv_2
XFILLER_167_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09173_ _09173_/A vssd1 vssd1 vccd1 vccd1 _10115_/A sky130_fd_sc_hd__buf_4
XANTENNA__11098__S0 _09447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13164__B2 _18621_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12396__A1_N _14584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14416__A1 _18516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12111__B _13608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10850_ _10850_/A _10850_/B vssd1 vssd1 vccd1 vccd1 _10850_/X sky130_fd_sc_hd__or2_1
XFILLER_44_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09509_ _09679_/A vssd1 vssd1 vccd1 vccd1 _10498_/A sky130_fd_sc_hd__clkbuf_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10781_ _10589_/A _10767_/X _10780_/X vssd1 vssd1 vccd1 vccd1 _10781_/X sky130_fd_sc_hd__a21bo_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14319__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12520_ _12520_/A vssd1 vssd1 vccd1 vccd1 _12751_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_12_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12451_ _19759_/Q _12451_/B vssd1 vssd1 vccd1 vccd1 _12451_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11402_ _12520_/A _11413_/A _12751_/D vssd1 vssd1 vccd1 vccd1 _12526_/A sky130_fd_sc_hd__nor3_4
X_15170_ _15170_/A vssd1 vssd1 vccd1 vccd1 _18660_/D sky130_fd_sc_hd__clkbuf_1
X_12382_ _12383_/A _14300_/B vssd1 vssd1 vccd1 vccd1 _12384_/A sky130_fd_sc_hd__and2_1
XFILLER_125_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14121_ _13966_/X _13968_/X _14121_/S vssd1 vssd1 vccd1 vccd1 _14121_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11333_ _11534_/B _11339_/B _11322_/D vssd1 vssd1 vccd1 vccd1 _11333_/X sky130_fd_sc_hd__or3b_2
XFILLER_21_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09148__A _09841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14052_ _18435_/Q _14050_/X _14209_/S vssd1 vssd1 vccd1 vccd1 _14053_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11264_ _10462_/A _11242_/Y _11132_/Y vssd1 vssd1 vccd1 vccd1 _11264_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_140_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13003_ _18314_/Q _13003_/B _13003_/C vssd1 vssd1 vccd1 vccd1 _13004_/C sky130_fd_sc_hd__and3_1
X_10215_ _10270_/A _10215_/B vssd1 vssd1 vccd1 vccd1 _10215_/X sky130_fd_sc_hd__or2_1
XANTENNA__15584__S _15584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17365__A _17376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18860_ _19543_/CLK _18860_/D vssd1 vssd1 vccd1 vccd1 _18860_/Q sky130_fd_sc_hd__dfxtp_1
X_11195_ _09317_/A _11185_/Y _11190_/X _11194_/Y _09394_/A vssd1 vssd1 vccd1 vccd1
+ _11195_/X sky130_fd_sc_hd__o311a_1
XFILLER_122_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17811_ _17811_/A vssd1 vssd1 vccd1 vccd1 _19707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10146_ _10127_/A _10145_/X _09621_/X vssd1 vssd1 vccd1 vccd1 _10146_/Y sky130_fd_sc_hd__o21ai_1
X_18791_ _19539_/CLK _18791_/D vssd1 vssd1 vccd1 vccd1 _18791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output143_A _11557_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17742_ _18483_/Q _17743_/B vssd1 vssd1 vccd1 vccd1 _17751_/C sky130_fd_sc_hd__or2_2
XFILLER_153_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14954_ _14954_/A vssd1 vssd1 vccd1 vccd1 _18606_/D sky130_fd_sc_hd__clkbuf_1
X_10077_ _09173_/A _10076_/X _09996_/A vssd1 vssd1 vccd1 vccd1 _10077_/X sky130_fd_sc_hd__a21o_1
XFILLER_130_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13905_ _14135_/A _13667_/X _13806_/A vssd1 vssd1 vccd1 vccd1 _13905_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17673_ _18471_/Q _17674_/B vssd1 vssd1 vccd1 vccd1 _17683_/C sky130_fd_sc_hd__or2_2
X_14885_ _18441_/Q _13305_/B _14992_/S vssd1 vssd1 vccd1 vccd1 _14885_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16709__A _16709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19412_ _19659_/CLK _19412_/D vssd1 vssd1 vccd1 vccd1 _19412_/Q sky130_fd_sc_hd__dfxtp_1
X_16624_ _16624_/A vssd1 vssd1 vccd1 vccd1 _19267_/D sky130_fd_sc_hd__clkbuf_1
X_13836_ _13881_/S _13836_/B vssd1 vssd1 vccd1 vccd1 _13836_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19343_ _19700_/CLK _19343_/D vssd1 vssd1 vccd1 vccd1 _19343_/Q sky130_fd_sc_hd__dfxtp_1
X_16555_ _16555_/A vssd1 vssd1 vccd1 vccd1 _19233_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13767_ _13618_/X _13636_/X _13768_/S vssd1 vssd1 vccd1 vccd1 _13767_/X sky130_fd_sc_hd__mux2_1
X_10979_ _12462_/A _11070_/A _12463_/A _11696_/A vssd1 vssd1 vccd1 vccd1 _10979_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_149_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15506_ _16761_/A vssd1 vssd1 vccd1 vccd1 _15506_/X sky130_fd_sc_hd__buf_2
X_19274_ _19628_/CLK _19274_/D vssd1 vssd1 vccd1 vccd1 _19274_/Q sky130_fd_sc_hd__dfxtp_1
X_12718_ _13426_/A _18631_/Q vssd1 vssd1 vccd1 vccd1 _12718_/Y sky130_fd_sc_hd__nand2_1
X_16486_ _16112_/X _19203_/Q _16486_/S vssd1 vssd1 vccd1 vccd1 _16487_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13698_ _13702_/A _13720_/B vssd1 vssd1 vccd1 vccd1 _13922_/B sky130_fd_sc_hd__or2_2
X_18225_ _18225_/A vssd1 vssd1 vccd1 vccd1 _18250_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15437_ _18762_/Q _15168_/X _15437_/S vssd1 vssd1 vccd1 vccd1 _15438_/A sky130_fd_sc_hd__mux2_1
X_12649_ _19780_/Q _12666_/B _12648_/X vssd1 vssd1 vccd1 vccd1 _14946_/B sky130_fd_sc_hd__o21a_2
XANTENNA__16444__A _16501_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18156_ _19839_/Q _19838_/Q _18156_/C vssd1 vssd1 vccd1 vccd1 _18158_/B sky130_fd_sc_hd__and3_1
XFILLER_157_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15368_ _15368_/A vssd1 vssd1 vccd1 vccd1 _18732_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09693__S0 _10257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11588__A _12458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17107_ _17107_/A vssd1 vssd1 vccd1 vccd1 _19453_/D sky130_fd_sc_hd__clkbuf_1
X_14319_ _14319_/A _14319_/B vssd1 vssd1 vccd1 vccd1 _14319_/Y sky130_fd_sc_hd__nor2_1
X_18087_ _18086_/B _18086_/C _19815_/Q vssd1 vssd1 vccd1 vccd1 _18088_/C sky130_fd_sc_hd__a21oi_1
XFILLER_144_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15299_ _15299_/A vssd1 vssd1 vccd1 vccd1 _18702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17038_ _17049_/A vssd1 vssd1 vccd1 vccd1 _17047_/S sky130_fd_sc_hd__buf_6
XFILLER_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_74_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09860_ _19622_/Q _19460_/Q _18906_/Q _18676_/Q _09911_/S _09841_/A vssd1 vssd1 vccd1
+ vccd1 _09861_/B sky130_fd_sc_hd__mux4_1
XFILLER_131_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10904__B1 _09625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09492__S _10511_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09791_ _18841_/Q _19395_/Q _19557_/Q _18809_/Q _09760_/X _09763_/X vssd1 vssd1 vccd1
+ vccd1 _09791_/X sky130_fd_sc_hd__mux4_2
XFILLER_113_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18989_ _19442_/CLK _18989_/D vssd1 vssd1 vccd1 vccd1 _18989_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09748__S1 _10186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15523__A _15590_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15071__A1 _13435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10667__A _10905_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13043__A _18085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09225_ _09225_/A vssd1 vssd1 vccd1 vccd1 _09459_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09156_ _10465_/S vssd1 vssd1 vccd1 vccd1 _09643_/S sky130_fd_sc_hd__buf_2
XFILLER_108_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10818__S0 _10982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12593__C1 _12592_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11498__A _18564_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09087_ _11314_/A vssd1 vssd1 vccd1 vccd1 _13570_/A sky130_fd_sc_hd__buf_4
XFILLER_135_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14885__A1 _13305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10046__S1 _10029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09987__S1 _09984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10000_ _09992_/A _09999_/X _09231_/A vssd1 vssd1 vccd1 vccd1 _10000_/X sky130_fd_sc_hd__o21a_1
XFILLER_153_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09989_ _09908_/A _09987_/X _09988_/X vssd1 vssd1 vccd1 vccd1 _09989_/X sky130_fd_sc_hd__o21a_1
XANTENNA__14637__B2 _14543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12648__B1 _13123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ _11953_/A _13620_/A vssd1 vssd1 vccd1 vccd1 _11952_/A sky130_fd_sc_hd__or2_1
XFILLER_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17124__S _17130_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10902_ _10895_/Y _10897_/Y _10899_/Y _10901_/Y _10846_/A vssd1 vssd1 vccd1 vccd1
+ _10902_/X sky130_fd_sc_hd__o221a_1
X_11882_ _11901_/A _11901_/C vssd1 vssd1 vccd1 vccd1 _11882_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_33_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14670_ _14670_/A vssd1 vssd1 vccd1 vccd1 _18576_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13621_ _14074_/B _12180_/A _13682_/S vssd1 vssd1 vccd1 vccd1 _13621_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17339__A0 _16771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10833_ _10825_/X _10828_/X _10830_/X _10832_/X _09244_/A vssd1 vssd1 vccd1 vccd1
+ _10833_/X sky130_fd_sc_hd__a221o_1
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09816__A1 _09819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12495__C _12495_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16340_ _16112_/X _19139_/Q _16340_/S vssd1 vssd1 vccd1 vccd1 _16341_/A sky130_fd_sc_hd__mux2_1
X_10764_ _10764_/A _10764_/B vssd1 vssd1 vccd1 vccd1 _10764_/Y sky130_fd_sc_hd__nor2_1
X_13552_ _13552_/A vssd1 vssd1 vccd1 vccd1 _18421_/D sky130_fd_sc_hd__clkbuf_1
X_12503_ _12503_/A _12503_/B vssd1 vssd1 vccd1 vccd1 _12503_/Y sky130_fd_sc_hd__nor2_1
X_13483_ _13483_/A vssd1 vssd1 vccd1 vccd1 _18400_/D sky130_fd_sc_hd__clkbuf_1
X_16271_ _16115_/X _19108_/Q _16279_/S vssd1 vssd1 vccd1 vccd1 _16272_/A sky130_fd_sc_hd__mux2_1
X_10695_ _10695_/A vssd1 vssd1 vccd1 vccd1 _11065_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18010_ _19788_/Q _18011_/C _18009_/Y vssd1 vssd1 vccd1 vccd1 _19788_/D sky130_fd_sc_hd__o21a_1
X_15222_ _15222_/A vssd1 vssd1 vccd1 vccd1 _18676_/D sky130_fd_sc_hd__clkbuf_1
X_12434_ _19758_/Q _12434_/B vssd1 vssd1 vccd1 vccd1 _12451_/B sky130_fd_sc_hd__nand2_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17794__S _17794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12365_ _19686_/Q _11989_/X _12364_/X _12193_/X vssd1 vssd1 vccd1 vccd1 _12365_/X
+ sky130_fd_sc_hd__o211a_1
X_15153_ _18655_/Q _15152_/X _15153_/S vssd1 vssd1 vccd1 vccd1 _15154_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15117__A2 _15116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14104_ _13750_/X _13952_/X _14103_/Y _13999_/S vssd1 vssd1 vccd1 vccd1 _14104_/X
+ sky130_fd_sc_hd__a211o_1
X_11316_ _11343_/C _11484_/B vssd1 vssd1 vccd1 vccd1 _11551_/B sky130_fd_sc_hd__and2_1
X_15084_ _18620_/Q _15083_/X _15087_/S vssd1 vssd1 vccd1 vccd1 _15085_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12296_ _11980_/X _12294_/X _12295_/X vssd1 vssd1 vccd1 vccd1 _12296_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18912_ _19628_/CLK _18912_/D vssd1 vssd1 vccd1 vccd1 _18912_/Q sky130_fd_sc_hd__dfxtp_1
X_14035_ _14035_/A vssd1 vssd1 vccd1 vccd1 _14035_/Y sky130_fd_sc_hd__inv_2
X_11247_ _11247_/A _11247_/B vssd1 vssd1 vccd1 vccd1 _11261_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__16203__S _16205_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09752__B1 _09625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16430__C _16919_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18843_ _19397_/CLK _18843_/D vssd1 vssd1 vccd1 vccd1 _18843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11178_ _11178_/A _11178_/B vssd1 vssd1 vccd1 vccd1 _11178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10129_ _18868_/Q _19326_/Q _10129_/S vssd1 vssd1 vccd1 vccd1 _10130_/A sky130_fd_sc_hd__mux2_1
X_18774_ _19295_/CLK _18774_/D vssd1 vssd1 vccd1 vccd1 _18774_/Q sky130_fd_sc_hd__dfxtp_1
X_15986_ _14833_/X _18992_/Q _15994_/S vssd1 vssd1 vccd1 vccd1 _15987_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17725_ _17713_/X _13334_/X _17724_/X vssd1 vssd1 vccd1 vccd1 _17725_/X sky130_fd_sc_hd__a21bo_1
X_14937_ input11/X _14901_/X _14904_/X vssd1 vssd1 vccd1 vccd1 _14937_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_36_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17034__S _17036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17656_ _18468_/Q _17656_/B vssd1 vssd1 vccd1 vccd1 _17657_/B sky130_fd_sc_hd__nand2_1
X_14868_ _14867_/X _18599_/Q _14880_/S vssd1 vssd1 vccd1 vccd1 _14869_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11862__B2 _11514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09341__A _10277_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16607_ _19259_/Q vssd1 vssd1 vccd1 vccd1 _16608_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_90_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13819_ _13899_/A vssd1 vssd1 vccd1 vccd1 _13819_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17587_ _17587_/A vssd1 vssd1 vccd1 vccd1 _19651_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13064__B1 _13063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14799_ _14825_/A vssd1 vssd1 vccd1 vccd1 _14980_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19326_ _19326_/CLK _19326_/D vssd1 vssd1 vccd1 vccd1 _19326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16538_ _16560_/A vssd1 vssd1 vccd1 vccd1 _16547_/S sky130_fd_sc_hd__buf_4
XANTENNA__11614__A1 _18562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09902__S1 _09783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13798__A _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10822__C1 _10821_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19257_ _19708_/CLK _19257_/D vssd1 vssd1 vccd1 vccd1 _19257_/Q sky130_fd_sc_hd__dfxtp_1
X_16469_ _16087_/X _19195_/Q _16475_/S vssd1 vssd1 vccd1 vccd1 _16470_/A sky130_fd_sc_hd__mux2_1
X_18208_ _19857_/Q _18214_/B vssd1 vssd1 vccd1 vccd1 _18210_/A sky130_fd_sc_hd__and2_1
XFILLER_164_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19188_ _19712_/CLK _19188_/D vssd1 vssd1 vccd1 vccd1 _19188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18139_ _18140_/B _18140_/C _19833_/Q vssd1 vssd1 vccd1 vccd1 _18141_/B sky130_fd_sc_hd__a21oi_1
XFILLER_156_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11111__A _11111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09912_ _09149_/A _09911_/X _09788_/A vssd1 vssd1 vccd1 vccd1 _09912_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_137_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16113__S _16113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10950__A _10950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11765__B _15255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09843_ _09843_/A _09843_/B vssd1 vssd1 vccd1 vccd1 _09843_/X sky130_fd_sc_hd__and2_1
XFILLER_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14619__A1 _11511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _10093_/A vssd1 vssd1 vccd1 vccd1 _09908_/A sky130_fd_sc_hd__clkbuf_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13980__B _13984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11066__C1 _10793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09208_ _09208_/A vssd1 vssd1 vccd1 vccd1 _09209_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_155_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10480_ _11102_/A _10480_/B vssd1 vssd1 vccd1 vccd1 _10480_/X sky130_fd_sc_hd__or2_1
XFILLER_6_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09139_ _09139_/A vssd1 vssd1 vccd1 vccd1 _10422_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10267__S1 _09145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ _13316_/A _12169_/C _11994_/A vssd1 vssd1 vccd1 vccd1 _12150_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11101_ _19610_/Q _19448_/Q _18894_/Q _18664_/Q _09449_/A _09538_/A vssd1 vssd1 vccd1
+ vccd1 _11102_/B sky130_fd_sc_hd__mux4_1
XANTENNA__17119__S _17119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10019__S1 _09979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15428__A _15485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ _12106_/A _12081_/B vssd1 vssd1 vccd1 vccd1 _12082_/B sky130_fd_sc_hd__or2_1
XFILLER_2_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16023__S _16027_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11032_ _19403_/Q _19179_/Q _19696_/Q _19147_/Q _10983_/S _10739_/A vssd1 vssd1 vccd1
+ vccd1 _11032_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16958__S _16964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10659__A1_N _18434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15840_ _15840_/A vssd1 vssd1 vccd1 vccd1 _18926_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19643_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__15283__A1 _15159_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _15793_/A vssd1 vssd1 vccd1 vccd1 _15780_/S sky130_fd_sc_hd__buf_4
XFILLER_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ _12983_/A _12983_/B _12983_/C vssd1 vssd1 vccd1 vccd1 _18308_/D sky130_fd_sc_hd__nor3_1
XFILLER_57_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _19617_/Q _16705_/X _17518_/S vssd1 vssd1 vccd1 vccd1 _17511_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14722_ _15077_/S vssd1 vssd1 vccd1 vccd1 _14762_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_73_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _19669_/Q _11959_/B vssd1 vssd1 vccd1 vccd1 _11934_/X sky130_fd_sc_hd__or2_1
X_18490_ _19468_/CLK _18490_/D vssd1 vssd1 vccd1 vccd1 _18490_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09161__A _10011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_22_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _17441_/A vssd1 vssd1 vccd1 vccd1 _19586_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14653_ _14555_/A _14648_/X _14649_/X input42/X vssd1 vssd1 vccd1 vccd1 _17777_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _14005_/B _11939_/B vssd1 vssd1 vccd1 vccd1 _11866_/B sky130_fd_sc_hd__nor2_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output106_A _09109_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13597__A1 _14176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13604_ _13604_/A vssd1 vssd1 vccd1 vccd1 _14155_/B sky130_fd_sc_hd__buf_2
X_17372_ _16819_/X _19556_/Q _17374_/S vssd1 vssd1 vccd1 vccd1 _17373_/A sky130_fd_sc_hd__mux2_1
X_10816_ _19247_/Q _19018_/Q _18949_/Q _19343_/Q _10982_/S _10969_/A vssd1 vssd1 vccd1
+ vccd1 _10816_/X sky130_fd_sc_hd__mux4_1
X_11796_ _19664_/Q _11795_/X _12191_/A vssd1 vssd1 vccd1 vccd1 _11796_/X sky130_fd_sc_hd__mux2_1
X_14584_ _14584_/A _14589_/B vssd1 vssd1 vccd1 vccd1 _14584_/X sky130_fd_sc_hd__or2_1
XFILLER_32_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19111_ _19657_/CLK _19111_/D vssd1 vssd1 vccd1 vccd1 _19111_/Q sky130_fd_sc_hd__dfxtp_1
X_16323_ _16087_/X _19131_/Q _16329_/S vssd1 vssd1 vccd1 vccd1 _16324_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13535_ _13535_/A vssd1 vssd1 vccd1 vccd1 _18417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10747_ _10750_/A _10746_/X _09224_/A vssd1 vssd1 vccd1 vccd1 _10747_/X sky130_fd_sc_hd__o21a_1
XFILLER_158_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19042_ _19657_/CLK _19042_/D vssd1 vssd1 vccd1 vccd1 _19042_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13411__A hold3/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16254_ _16254_/A vssd1 vssd1 vccd1 vccd1 _19100_/D sky130_fd_sc_hd__clkbuf_1
X_13466_ _13512_/S vssd1 vssd1 vccd1 vccd1 _13475_/S sky130_fd_sc_hd__clkbuf_4
X_10678_ _11027_/S vssd1 vssd1 vccd1 vccd1 _10860_/S sky130_fd_sc_hd__buf_2
XANTENNA__09648__S0 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15205_ _18671_/Q _15203_/X _15217_/S vssd1 vssd1 vccd1 vccd1 _15206_/A sky130_fd_sc_hd__mux2_1
X_12417_ _19757_/Q _11705_/X _12413_/X _12416_/Y vssd1 vssd1 vccd1 vccd1 _17909_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_127_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16185_ _16196_/A vssd1 vssd1 vccd1 vccd1 _16194_/S sky130_fd_sc_hd__buf_4
XANTENNA__14941__S _14941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17818__A _17840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13397_ _19788_/Q _13123_/X _13393_/X _13396_/X vssd1 vssd1 vccd1 vccd1 _13398_/B
+ sky130_fd_sc_hd__a211o_2
XANTENNA__16722__A _16722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15136_ _16138_/A _16212_/B _15960_/C vssd1 vssd1 vccd1 vccd1 _16503_/A sky130_fd_sc_hd__or3_4
X_12348_ _12348_/A vssd1 vssd1 vccd1 vccd1 _13712_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11866__A _11970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ _13567_/A _14241_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _12280_/B sky130_fd_sc_hd__o21ai_1
X_15067_ _15066_/X _18616_/Q _15077_/S vssd1 vssd1 vccd1 vccd1 _15068_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14018_ _14018_/A vssd1 vssd1 vccd1 vccd1 _14018_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17799__A0 _15159_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10335__A1 _09616_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15772__S _15780_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18826_ _19639_/CLK _18826_/D vssd1 vssd1 vccd1 vccd1 _18826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18757_ _19698_/CLK _18757_/D vssd1 vssd1 vccd1 vccd1 _18757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15969_ _15969_/A vssd1 vssd1 vccd1 vccd1 _18984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17708_ _17708_/A vssd1 vssd1 vccd1 vccd1 _17708_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09490_ _10788_/S vssd1 vssd1 vccd1 vccd1 _10500_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18688_ _19791_/CLK _18688_/D vssd1 vssd1 vccd1 vccd1 _18688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13305__B _13305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17639_ _18465_/Q _17640_/B vssd1 vssd1 vccd1 vccd1 _17649_/C sky130_fd_sc_hd__or2_2
XFILLER_24_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09887__S0 _09809_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19309_ _19691_/CLK _19309_/D vssd1 vssd1 vccd1 vccd1 _19309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10497__S1 _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12260__A1 _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11771__B1 _11997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13467__S _13475_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11776__A _11776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13512__A1 _13437_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09246__A _09246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10326__A1 _19194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09811__S0 _09809_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09826_ _09826_/A _09826_/B vssd1 vssd1 vccd1 vccd1 _09826_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17463__A _17463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10421__S1 _09142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09757_ _10257_/S vssd1 vssd1 vccd1 vccd1 _10094_/A sky130_fd_sc_hd__buf_2
XFILLER_74_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _09688_/A _12501_/A vssd1 vssd1 vccd1 vccd1 _09755_/A sky130_fd_sc_hd__nor2_1
XANTENNA__15017__A1 _18452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17402__S _17402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11070_/A _18492_/Q _11840_/A vssd1 vssd1 vccd1 vccd1 _13665_/A sky130_fd_sc_hd__mux2_4
XFILLER_30_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10601_ _12474_/B _10601_/B vssd1 vssd1 vccd1 vccd1 _10601_/X sky130_fd_sc_hd__and2b_1
XFILLER_167_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16517__A1 _15506_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11581_ _11579_/Y _11580_/X _18574_/Q _11575_/Y vssd1 vssd1 vccd1 vccd1 _11581_/Y
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__10488__S1 _09483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13320_ _12634_/B _13311_/X _13319_/X _13317_/X vssd1 vssd1 vccd1 vccd1 _18369_/D
+ sky130_fd_sc_hd__o211a_1
X_10532_ _09549_/A _10531_/X _09210_/A vssd1 vssd1 vccd1 vccd1 _10532_/X sky130_fd_sc_hd__o21a_1
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15857__S _15863_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13251_ _13251_/A vssd1 vssd1 vccd1 vccd1 _13251_/X sky130_fd_sc_hd__clkbuf_2
X_10463_ _19254_/Q _19025_/Q _18956_/Q _19350_/Q _09631_/A _10368_/A vssd1 vssd1 vccd1
+ vccd1 _10464_/B sky130_fd_sc_hd__mux4_1
XFILLER_6_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12202_ _18575_/Q _11966_/B _12173_/Y vssd1 vssd1 vccd1 vccd1 _12202_/X sky130_fd_sc_hd__a21o_1
X_13182_ _13121_/X _13171_/Y _13181_/X _13135_/X _18623_/Q vssd1 vssd1 vccd1 vccd1
+ _13182_/X sky130_fd_sc_hd__a32o_4
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input67_A io_irq_m1_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10394_ _10442_/A _10394_/B vssd1 vssd1 vccd1 vccd1 _10394_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_142_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19467_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_151_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12133_ _14178_/B _12133_/B vssd1 vssd1 vccd1 vccd1 _12137_/A sky130_fd_sc_hd__xnor2_1
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990_ _19782_/Q _17990_/B vssd1 vssd1 vccd1 vccd1 _17997_/C sky130_fd_sc_hd__and2_1
XFILLER_97_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16941_ _16941_/A vssd1 vssd1 vccd1 vccd1 _19379_/D sky130_fd_sc_hd__clkbuf_1
X_12064_ _12064_/A _12064_/B vssd1 vssd1 vccd1 vccd1 _12066_/A sky130_fd_sc_hd__nor2_2
XANTENNA__09156__A _10465_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10317__A1 _10080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11015_ _19630_/Q _19047_/Q _19084_/Q _18690_/Q _09336_/A _10940_/X vssd1 vssd1 vccd1
+ vccd1 _11016_/B sky130_fd_sc_hd__mux4_2
X_19660_ _19660_/CLK _19660_/D vssd1 vssd1 vccd1 vccd1 _19660_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_157_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19601_/CLK sky130_fd_sc_hd__clkbuf_16
X_16872_ _19349_/Q _16673_/X _16880_/S vssd1 vssd1 vccd1 vccd1 _16873_/A sky130_fd_sc_hd__mux2_1
X_18611_ _19554_/CLK _18611_/D vssd1 vssd1 vccd1 vccd1 _18611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15823_ _15823_/A vssd1 vssd1 vccd1 vccd1 _18918_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19591_ _19591_/CLK _19591_/D vssd1 vssd1 vccd1 vccd1 _19591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18542_ _19481_/CLK _18542_/D vssd1 vssd1 vccd1 vccd1 _18542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _14792_/X _18888_/Q _15758_/S vssd1 vssd1 vccd1 vccd1 _15755_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12966_ _14673_/A vssd1 vssd1 vccd1 vccd1 _14638_/A sky130_fd_sc_hd__buf_4
XFILLER_80_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10176__S0 _09721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _11046_/A _13134_/B _14922_/S vssd1 vssd1 vccd1 vccd1 _14705_/X sky130_fd_sc_hd__mux2_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _11918_/A _13622_/A vssd1 vssd1 vccd1 vccd1 _11919_/A sky130_fd_sc_hd__nand2_1
X_18473_ _19079_/CLK _18473_/D vssd1 vssd1 vccd1 vccd1 _18473_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15685_ _15685_/A vssd1 vssd1 vccd1 vccd1 _18857_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12897_ _12897_/A _12897_/B vssd1 vssd1 vccd1 vccd1 _12897_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17953__B1 _19769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17424_ _16790_/X _19579_/Q _17424_/S vssd1 vssd1 vccd1 vccd1 _17425_/A sky130_fd_sc_hd__mux2_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _14636_/A vssd1 vssd1 vccd1 vccd1 _18565_/D sky130_fd_sc_hd__clkbuf_1
X_11848_ _11849_/A _12095_/B _19735_/Q vssd1 vssd1 vccd1 vccd1 _11851_/A sky130_fd_sc_hd__a21oi_1
XFILLER_33_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15340__B _17391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17355_ _16793_/X _19548_/Q _17363_/S vssd1 vssd1 vccd1 vccd1 _17356_/A sky130_fd_sc_hd__mux2_1
X_14567_ _12540_/A _14564_/X _14566_/X _14560_/X vssd1 vssd1 vccd1 vccd1 _18543_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17705__A0 _19677_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16508__A1 _15494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11779_ _11779_/A vssd1 vssd1 vccd1 vccd1 _11779_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16306_ _16306_/A vssd1 vssd1 vccd1 vccd1 _19123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11450__C1 _11720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13518_ _18415_/Q _12731_/A _14526_/B _14431_/C _13542_/A vssd1 vssd1 vccd1 vccd1
+ _18415_/D sky130_fd_sc_hd__o221a_1
XANTENNA__13990__A1 _18432_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17286_ _17286_/A vssd1 vssd1 vccd1 vccd1 _19517_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17181__A1 _12727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14498_ _18519_/Q _19757_/Q _14498_/S vssd1 vssd1 vccd1 vccd1 _14499_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19025_ _19610_/CLK _19025_/D vssd1 vssd1 vccd1 vccd1 _19025_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15767__S _15769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16237_ _16283_/S vssd1 vssd1 vccd1 vccd1 _16246_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__17548__A _17605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13449_ _18385_/Q _13165_/Y _13453_/S vssd1 vssd1 vccd1 vccd1 _13450_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16168_ _16074_/X _19058_/Q _16172_/S vssd1 vssd1 vccd1 vccd1 _16169_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18130__B1 _19830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11753__B1 _19732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15119_ _18639_/Q _15116_/X _15118_/X _10098_/X vssd1 vssd1 vccd1 vccd1 _18639_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16099_ _16809_/A vssd1 vssd1 vccd1 vccd1 _16099_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15495__A1 _15494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19858_ _19858_/CLK _19858_/D vssd1 vssd1 vccd1 vccd1 _19858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09611_ _19530_/Q _19144_/Q _19594_/Q _18750_/Q _10131_/S _09610_/X vssd1 vssd1 vccd1
+ vccd1 _09612_/B sky130_fd_sc_hd__mux4_1
X_18809_ _19557_/CLK _18809_/D vssd1 vssd1 vccd1 vccd1 _18809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19789_ _19790_/CLK _19789_/D vssd1 vssd1 vccd1 vccd1 _19789_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16995__A1 _16639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09542_ _09542_/A vssd1 vssd1 vccd1 vccd1 _09978_/A sky130_fd_sc_hd__buf_4
XFILLER_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09473_ _10895_/A vssd1 vssd1 vccd1 vccd1 _10764_/A sky130_fd_sc_hd__buf_2
XFILLER_52_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10675__A _10875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10890__S1 _09512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__S _09675_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_74_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19810_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_133_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09809_ _09872_/S vssd1 vssd1 vccd1 vccd1 _09809_/X sky130_fd_sc_hd__buf_4
XANTENNA__09704__A _09704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11953__B _13620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_89_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _18329_/CLK sky130_fd_sc_hd__clkbuf_16
X_12820_ _12821_/B _12821_/C _18256_/Q vssd1 vssd1 vccd1 vccd1 _12822_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10158__S0 _10256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _14562_/A _12751_/B _12751_/C _12751_/D vssd1 vssd1 vccd1 vccd1 _12752_/A
+ sky130_fd_sc_hd__nor4_4
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17132__S _17134_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11702_ _11703_/B _11702_/B vssd1 vssd1 vccd1 vccd1 _11746_/B sky130_fd_sc_hd__and2b_2
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19624_/CLK sky130_fd_sc_hd__clkbuf_16
X_15470_ _18777_/Q _15216_/X _15470_/S vssd1 vssd1 vccd1 vccd1 _15471_/A sky130_fd_sc_hd__mux2_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _18306_/Q _12663_/X _12681_/X vssd1 vssd1 vccd1 vccd1 _12683_/B sky130_fd_sc_hd__a21oi_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14213__A2 _13623_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _18486_/Q _18518_/Q _14424_/S vssd1 vssd1 vccd1 vccd1 _14422_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _13625_/A _13789_/A _11940_/A vssd1 vssd1 vccd1 vccd1 _11648_/A sky130_fd_sc_hd__o21ai_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16971__S _16975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17140_ _17245_/S vssd1 vssd1 vccd1 vccd1 _17155_/S sky130_fd_sc_hd__buf_2
XFILLER_24_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14352_ _14765_/A _18494_/Q _14352_/S vssd1 vssd1 vccd1 vccd1 _14353_/A sky130_fd_sc_hd__mux2_1
X_11564_ _11564_/A _11575_/B vssd1 vssd1 vccd1 vccd1 _11565_/C sky130_fd_sc_hd__nor2_1
XANTENNA__11983__B1 _17878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13303_ _19674_/Q _12737_/X _13301_/X _13302_/X vssd1 vssd1 vccd1 vccd1 _13303_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_128_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_27_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19616_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15587__S _15590_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17071_ _16752_/X _19437_/Q _17075_/S vssd1 vssd1 vccd1 vccd1 _17072_/A sky130_fd_sc_hd__mux2_1
X_10515_ _18763_/Q _18992_/Q _18923_/Q _19221_/Q _10579_/S _10651_/A vssd1 vssd1 vccd1
+ vccd1 _10516_/B sky130_fd_sc_hd__mux4_1
XFILLER_144_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14283_ _14283_/A vssd1 vssd1 vccd1 vccd1 _18452_/D sky130_fd_sc_hd__clkbuf_1
X_11495_ _11511_/A _11495_/B vssd1 vssd1 vccd1 vccd1 _11664_/C sky130_fd_sc_hd__or2_1
XFILLER_109_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16022_ _16022_/A vssd1 vssd1 vccd1 vccd1 _19008_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09585__S _10125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13234_ _13248_/A _18628_/Q vssd1 vssd1 vccd1 vccd1 _13234_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10446_ _19255_/Q _19026_/Q _18957_/Q _19351_/Q _11112_/S _10384_/X vssd1 vssd1 vccd1
+ vccd1 _10447_/B sky130_fd_sc_hd__mux4_1
XFILLER_137_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13165_ _15254_/B vssd1 vssd1 vccd1 vccd1 _13165_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10002__A3 _10001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10377_ _10379_/A _10376_/X _09434_/X vssd1 vssd1 vccd1 vccd1 _10377_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12305__A _14265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12116_ _12116_/A vssd1 vssd1 vccd1 vccd1 _12116_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17973_ _19776_/Q _17973_/B vssd1 vssd1 vccd1 vccd1 _17979_/C sky130_fd_sc_hd__and2_1
XFILLER_124_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13096_ _17892_/A vssd1 vssd1 vccd1 vccd1 _17781_/A sky130_fd_sc_hd__buf_4
XANTENNA__18199__A _18199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12047_ _19673_/Q _11563_/X _17204_/A vssd1 vssd1 vccd1 vccd1 _12047_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__17307__S _17313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15616__A _15662_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16924_ _16924_/A vssd1 vssd1 vccd1 vccd1 _19371_/D sky130_fd_sc_hd__clkbuf_1
X_19712_ _19712_/CLK _19712_/D vssd1 vssd1 vccd1 vccd1 _19712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16855_ _16855_/A vssd1 vssd1 vccd1 vccd1 _19341_/D sky130_fd_sc_hd__clkbuf_1
X_19643_ _19643_/CLK _19643_/D vssd1 vssd1 vccd1 vccd1 _19643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15806_ _15076_/X _18912_/Q _15806_/S vssd1 vssd1 vccd1 vccd1 _15807_/A sky130_fd_sc_hd__mux2_1
X_19574_ _19726_/CLK _19574_/D vssd1 vssd1 vccd1 vccd1 _19574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16786_ _16786_/A vssd1 vssd1 vccd1 vccd1 _19319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13998_ _13816_/A _13996_/X _14135_/B _13838_/A vssd1 vssd1 vccd1 vccd1 _13998_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18525_ _19733_/CLK _18525_/D vssd1 vssd1 vccd1 vccd1 _18525_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15737_ _15793_/A vssd1 vssd1 vccd1 vccd1 _15806_/S sky130_fd_sc_hd__buf_6
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12949_ _18293_/Q _12952_/C _12948_/X vssd1 vssd1 vccd1 vccd1 _12949_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18456_ _19078_/CLK _18456_/D vssd1 vssd1 vccd1 vccd1 _18456_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_61_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15668_ _15668_/A vssd1 vssd1 vccd1 vccd1 _18849_/D sky130_fd_sc_hd__clkbuf_1
X_17407_ _16765_/X _19571_/Q _17413_/S vssd1 vssd1 vccd1 vccd1 _17408_/A sky130_fd_sc_hd__mux2_1
X_14619_ _11511_/A _14613_/X _14603_/X input63/X vssd1 vssd1 vccd1 vccd1 _14620_/B
+ sky130_fd_sc_hd__a22o_1
X_18387_ _19780_/CLK _18387_/D vssd1 vssd1 vccd1 vccd1 _18387_/Q sky130_fd_sc_hd__dfxtp_1
X_15599_ _18819_/Q _15497_/X _15603_/S vssd1 vssd1 vccd1 vccd1 _15600_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17338_ _17338_/A vssd1 vssd1 vccd1 vccd1 _19540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17154__A1 _13182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11974__A0 _10461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17269_ _19510_/Q _16670_/X _17269_/S vssd1 vssd1 vccd1 vccd1 _17270_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10872__S1 _10365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19008_ _19722_/CLK _19008_/D vssd1 vssd1 vccd1 vccd1 _19008_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_144_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12215__A _19747_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09524__A _10395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11773__B _15095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13100__C1 _14612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09525_ _10387_/S vssd1 vssd1 vccd1 vccd1 _10242_/S sky130_fd_sc_hd__buf_6
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13480__S _13486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_69_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09456_ _10622_/A vssd1 vssd1 vccd1 vccd1 _10574_/A sky130_fd_sc_hd__clkbuf_2
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09387_ _09814_/A _09386_/X _09320_/X vssd1 vssd1 vccd1 vccd1 _09387_/X sky130_fd_sc_hd__o21a_1
XFILLER_101_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16791__S _16791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10312__S0 _09701_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10300_ _10300_/A _10300_/B vssd1 vssd1 vccd1 vccd1 _11235_/A sky130_fd_sc_hd__nor2_1
XFILLER_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11280_ _11472_/A _11471_/A vssd1 vssd1 vccd1 vccd1 _11501_/B sky130_fd_sc_hd__nor2_2
XFILLER_118_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11717__B1 _11720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14324__B _14324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10231_ _10245_/A vssd1 vssd1 vccd1 vccd1 _11111_/A sky130_fd_sc_hd__buf_4
XFILLER_134_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10162_ _19519_/Q _19133_/Q _19583_/Q _18739_/Q _10200_/S _09146_/A vssd1 vssd1 vccd1
+ vccd1 _10163_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10093_ _10093_/A _10093_/B vssd1 vssd1 vccd1 vccd1 _10093_/X sky130_fd_sc_hd__or2_1
XANTENNA__16031__S _16031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14970_ _18448_/Q _13345_/B _14981_/S vssd1 vssd1 vccd1 vccd1 _14970_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13921_ _14130_/A _14293_/B vssd1 vssd1 vccd1 vccd1 _13931_/B sky130_fd_sc_hd__nor2_1
XFILLER_47_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12693__A1 _13104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11040__S1 _10969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12693__B2 _12692_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15870__S _15874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16640_ _16744_/A _16847_/B vssd1 vssd1 vccd1 vccd1 _16722_/A sky130_fd_sc_hd__nor2_4
X_13852_ _13993_/A vssd1 vssd1 vccd1 vccd1 _13966_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_75_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10299__B _12485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12803_ _12808_/B _18250_/B _12802_/X vssd1 vssd1 vccd1 vccd1 _12803_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13642__A0 _13671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16571_ _19241_/Q _15586_/X _16573_/S vssd1 vssd1 vccd1 vccd1 _16572_/A sky130_fd_sc_hd__mux2_1
X_13783_ _14102_/A _13783_/B vssd1 vssd1 vccd1 vccd1 _14097_/A sky130_fd_sc_hd__nor2_1
X_10995_ _18818_/Q _19372_/Q _19534_/Q _18786_/Q _10959_/X _10960_/X vssd1 vssd1 vccd1
+ vccd1 _10996_/B sky130_fd_sc_hd__mux4_1
X_18310_ _19795_/CLK _18310_/D vssd1 vssd1 vccd1 vccd1 _18310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15171__A _16673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15522_ _16777_/A vssd1 vssd1 vccd1 vccd1 _15522_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ _12734_/A _12751_/B _12751_/C _12751_/D vssd1 vssd1 vccd1 vccd1 _12735_/A
+ sky130_fd_sc_hd__nor4_4
X_19290_ _19612_/CLK _19290_/D vssd1 vssd1 vccd1 vccd1 _19290_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _18249_/A _18241_/B _18241_/C vssd1 vssd1 vccd1 vccd1 _19868_/D sky130_fd_sc_hd__nor3_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17797__S _17805_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14198__A1 _18445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13403__B hold3/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _18769_/Q _15191_/X _15459_/S vssd1 vssd1 vccd1 vccd1 _15454_/A sky130_fd_sc_hd__mux2_1
X_12665_ _12665_/A vssd1 vssd1 vccd1 vccd1 _12665_/X sky130_fd_sc_hd__buf_2
XFILLER_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14404_ _17728_/A _18512_/Q _14410_/S vssd1 vssd1 vccd1 vccd1 _14405_/A sky130_fd_sc_hd__mux2_1
X_18172_ _19844_/Q _18175_/C _18171_/Y vssd1 vssd1 vccd1 vccd1 _19844_/D sky130_fd_sc_hd__o21a_1
X_11616_ _11688_/C vssd1 vssd1 vccd1 vccd1 _13769_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__17136__A1 _13136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15384_ _18740_/Q _15200_/X _15384_/S vssd1 vssd1 vccd1 vccd1 _15385_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12596_ _13306_/A vssd1 vssd1 vccd1 vccd1 _12596_/X sky130_fd_sc_hd__clkbuf_2
X_17123_ _17123_/A vssd1 vssd1 vccd1 vccd1 _19460_/D sky130_fd_sc_hd__clkbuf_1
X_14335_ _14331_/Y _13806_/X _14334_/X _12447_/B _14000_/X vssd1 vssd1 vccd1 vccd1
+ _14335_/X sky130_fd_sc_hd__o2111a_1
XFILLER_156_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11547_ _15060_/B vssd1 vssd1 vccd1 vccd1 _15071_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17054_ _19430_/Q _16728_/X _17058_/S vssd1 vssd1 vccd1 vccd1 _17055_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output98_A _11704_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14266_ _14078_/A _14261_/Y _14265_/Y vssd1 vssd1 vccd1 vccd1 _14266_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11478_ _11478_/A _11598_/B vssd1 vssd1 vccd1 vccd1 _13520_/A sky130_fd_sc_hd__or2_1
X_16005_ _14940_/X _19001_/Q _16005_/S vssd1 vssd1 vccd1 vccd1 _16006_/A sky130_fd_sc_hd__mux2_1
X_13217_ _13297_/A vssd1 vssd1 vccd1 vccd1 _13217_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14370__A1 _18500_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10429_ _19641_/Q _19058_/Q _19095_/Q _18701_/Q _09632_/A _10368_/X vssd1 vssd1 vccd1
+ vccd1 _10429_/X sky130_fd_sc_hd__mux4_1
X_14197_ _12163_/Y _14070_/X _14196_/X _14099_/X vssd1 vssd1 vccd1 vccd1 _14197_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_124_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13148_ _18620_/Q _13148_/B vssd1 vssd1 vccd1 vccd1 _13148_/X sky130_fd_sc_hd__or2_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10931__B2 _18428_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13079_ _18342_/Q _12568_/X _12642_/A _13215_/A vssd1 vssd1 vccd1 vccd1 _13079_/X
+ sky130_fd_sc_hd__a22o_1
X_17956_ _17999_/A vssd1 vssd1 vccd1 vccd1 _17991_/A sky130_fd_sc_hd__clkbuf_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09344__A _09344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16907_ _19365_/Q _16725_/X _16913_/S vssd1 vssd1 vccd1 vccd1 _16908_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17887_ _12095_/A _17886_/X _12102_/X _14585_/X vssd1 vssd1 vccd1 vccd1 _19744_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12684__A1 _12766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11031__S1 _10960_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16876__S _16880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15780__S _15780_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19626_ _19626_/CLK _19626_/D vssd1 vssd1 vccd1 vccd1 _19626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16838_ _16838_/A vssd1 vssd1 vccd1 vccd1 _16838_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19557_ _19557_/CLK _19557_/D vssd1 vssd1 vccd1 vccd1 _19557_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13633__A0 _11784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16769_ _16768_/X _19314_/Q _16775_/S vssd1 vssd1 vccd1 vccd1 _16770_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09837__C1 _09395_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09310_ _18980_/Q vssd1 vssd1 vccd1 vccd1 _10728_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_70_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18508_ _18510_/CLK _18508_/D vssd1 vssd1 vccd1 vccd1 _18508_/Q sky130_fd_sc_hd__dfxtp_1
X_19488_ _19488_/CLK _19488_/D vssd1 vssd1 vccd1 vccd1 _19488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09241_ _09237_/A _09238_/X _09240_/X _09231_/X vssd1 vssd1 vccd1 vccd1 _09241_/X
+ sky130_fd_sc_hd__o211a_1
X_18439_ _19078_/CLK _18439_/D vssd1 vssd1 vccd1 vccd1 _18439_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13397__C1 _13396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09172_ _09172_/A vssd1 vssd1 vccd1 vccd1 _09173_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16640__A _16744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13475__S _13475_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11784__A _11784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13624__A0 _14057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09508_ _10638_/A vssd1 vssd1 vccd1 vccd1 _09679_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _10846_/A _10780_/B _10780_/C vssd1 vssd1 vccd1 vccd1 _10780_/X sky130_fd_sc_hd__or3_1
XFILLER_24_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _09629_/A vssd1 vssd1 vccd1 vccd1 _10540_/S sky130_fd_sc_hd__buf_2
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12450_ _12450_/A _12450_/B vssd1 vssd1 vccd1 vccd1 _12450_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_166_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11401_ _11401_/A vssd1 vssd1 vccd1 vccd1 _12751_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__11959__A _19670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10863__A _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12381_ _12381_/A vssd1 vssd1 vccd1 vccd1 _14300_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_153_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14120_ _14120_/A vssd1 vssd1 vccd1 vccd1 _14120_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_165_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11332_ _13526_/B _11344_/A _11519_/B vssd1 vssd1 vccd1 vccd1 _11585_/D sky130_fd_sc_hd__or3_2
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13155__A2 _13235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14051_ _15093_/S vssd1 vssd1 vccd1 vccd1 _14209_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_106_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11263_ _11263_/A _11263_/B vssd1 vssd1 vccd1 vccd1 _11263_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13002_ _13003_/B _13003_/C _18314_/Q vssd1 vssd1 vccd1 vccd1 _13004_/B sky130_fd_sc_hd__a21oi_1
XFILLER_122_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10214_ _19614_/Q _19452_/Q _18898_/Q _18668_/Q _09545_/S _09697_/A vssd1 vssd1 vccd1
+ vccd1 _10215_/B sky130_fd_sc_hd__mux4_1
XFILLER_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11194_ _11180_/A _11191_/X _11193_/X vssd1 vssd1 vccd1 vccd1 _11194_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_122_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10145_ _19616_/Q _19454_/Q _18900_/Q _18670_/Q _10125_/X _09595_/A vssd1 vssd1 vccd1
+ vccd1 _10145_/X sky130_fd_sc_hd__mux4_1
X_17810_ _15175_/X _19707_/Q _17816_/S vssd1 vssd1 vccd1 vccd1 _17811_/A sky130_fd_sc_hd__mux2_1
X_18790_ _19540_/CLK _18790_/D vssd1 vssd1 vccd1 vccd1 _18790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17741_ _19683_/Q _17708_/X _17739_/Y _17740_/X vssd1 vssd1 vccd1 vccd1 _19683_/D
+ sky130_fd_sc_hd__o22a_1
X_14953_ _14951_/X _18606_/Q _14997_/S vssd1 vssd1 vccd1 vccd1 _14954_/A sky130_fd_sc_hd__mux2_1
X_10076_ _18869_/Q _19327_/Q _10076_/S vssd1 vssd1 vccd1 vccd1 _10076_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13904_ _13753_/X _13667_/X _14323_/A vssd1 vssd1 vccd1 vccd1 _13904_/Y sky130_fd_sc_hd__a21oi_1
X_17672_ _17672_/A vssd1 vssd1 vccd1 vccd1 _19671_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10103__A _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14884_ _14883_/A _14894_/C _14815_/A vssd1 vssd1 vccd1 vccd1 _14884_/X sky130_fd_sc_hd__o21a_1
XFILLER_48_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16623_ _19267_/Q vssd1 vssd1 vccd1 vccd1 _16624_/A sky130_fd_sc_hd__clkbuf_1
X_19411_ _19571_/CLK _19411_/D vssd1 vssd1 vccd1 vccd1 _19411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13835_ _13663_/X _13669_/X _13877_/S vssd1 vssd1 vccd1 vccd1 _13836_/B sky130_fd_sc_hd__mux2_1
XFILLER_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12418__B2 _12504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16554_ _19233_/Q _15561_/X _16558_/S vssd1 vssd1 vccd1 vccd1 _16555_/A sky130_fd_sc_hd__mux2_1
X_19342_ _19568_/CLK _19342_/D vssd1 vssd1 vccd1 vccd1 _19342_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13766_ _13764_/X _13765_/X _13769_/S vssd1 vssd1 vccd1 vccd1 _13766_/X sky130_fd_sc_hd__mux2_1
X_10978_ _18429_/Q _09280_/A _10857_/X _10977_/X vssd1 vssd1 vccd1 vccd1 _11696_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_16_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15505_ _15505_/A vssd1 vssd1 vccd1 vccd1 _18789_/D sky130_fd_sc_hd__clkbuf_1
X_12717_ _17774_/A _18301_/Q _13090_/S _12716_/X vssd1 vssd1 vccd1 vccd1 _18301_/D
+ sky130_fd_sc_hd__o31a_1
X_19273_ _19713_/CLK _19273_/D vssd1 vssd1 vccd1 vccd1 _19273_/Q sky130_fd_sc_hd__dfxtp_1
X_16485_ _16485_/A vssd1 vssd1 vccd1 vccd1 _19202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13697_ _13720_/A _13785_/A vssd1 vssd1 vccd1 vccd1 _13870_/B sky130_fd_sc_hd__or2_1
XANTENNA__16725__A _16725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18224_ _19862_/Q _18221_/A _18223_/Y vssd1 vssd1 vccd1 vccd1 _19862_/D sky130_fd_sc_hd__o21a_1
X_15436_ _15436_/A vssd1 vssd1 vccd1 vccd1 _18761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12648_ _18287_/Q _12638_/X _13123_/A _12647_/X vssd1 vssd1 vccd1 vccd1 _12648_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18155_ _19838_/Q _18156_/C _19839_/Q vssd1 vssd1 vccd1 vccd1 _18157_/B sky130_fd_sc_hd__a21oi_1
XFILLER_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15367_ _18732_/Q _15175_/X _15373_/S vssd1 vssd1 vccd1 vccd1 _15368_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12579_ _13415_/A _18636_/Q vssd1 vssd1 vccd1 vccd1 _12579_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09693__S1 _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17106_ _16803_/X _19453_/Q _17108_/S vssd1 vssd1 vccd1 vccd1 _17107_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14318_ _09626_/Y _13873_/X _14317_/X vssd1 vssd1 vccd1 vccd1 _18455_/D sky130_fd_sc_hd__a21oi_1
XFILLER_172_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18086_ _19815_/Q _18086_/B _18086_/C vssd1 vssd1 vccd1 vccd1 _18088_/B sky130_fd_sc_hd__and3_1
XFILLER_144_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15298_ _18702_/Q _15181_/X _15300_/S vssd1 vssd1 vccd1 vccd1 _15299_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17037_ _17037_/A vssd1 vssd1 vccd1 vccd1 _19422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14249_ _12280_/A _14253_/A vssd1 vssd1 vccd1 vccd1 _14249_/X sky130_fd_sc_hd__and2b_1
XFILLER_125_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_17_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _09861_/A _09790_/B vssd1 vssd1 vccd1 vccd1 _09790_/X sky130_fd_sc_hd__or2_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _19539_/CLK _18988_/D vssd1 vssd1 vccd1 vccd1 _18988_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _19764_/Q _17935_/C _17938_/Y vssd1 vssd1 vccd1 vccd1 _19764_/D sky130_fd_sc_hd__o21a_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11109__A _11119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10763__S0 _10650_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09802__A _10033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13606__A0 _14138_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19609_ _19609_/CLK _19609_/D vssd1 vssd1 vccd1 vccd1 _19609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09224_ _09224_/A vssd1 vssd1 vccd1 vccd1 _09225_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_148_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09155_ _10466_/S vssd1 vssd1 vccd1 vccd1 _10465_/S sky130_fd_sc_hd__buf_4
XFILLER_147_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10818__S1 _10969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10683__A _10875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09249__A _09249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11498__B _18562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09086_ _09107_/A _11358_/B _12471_/B vssd1 vssd1 vccd1 vccd1 _11314_/A sky130_fd_sc_hd__nor3_2
XFILLER_174_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13137__A2 _13136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09988_ _09988_/A vssd1 vssd1 vccd1 vccd1 _09988_/X sky130_fd_sc_hd__buf_2
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12648__A1 _18287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13218__B _18627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17405__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__B1 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950_ _11082_/B _12060_/A _11949_/X vssd1 vssd1 vccd1 vccd1 _13620_/A sky130_fd_sc_hd__o21ai_4
XFILLER_83_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10754__S0 _09152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09712__A _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ _10895_/A _10900_/X _10793_/X vssd1 vssd1 vccd1 vccd1 _10901_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11881_ _19736_/Q vssd1 vssd1 vccd1 vccd1 _11901_/A sky130_fd_sc_hd__buf_4
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13620_ _13620_/A vssd1 vssd1 vccd1 vccd1 _14074_/B sky130_fd_sc_hd__inv_2
X_10832_ _10866_/A _10831_/X _10821_/X vssd1 vssd1 vccd1 vccd1 _10832_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13551_ _13560_/A _13551_/B vssd1 vssd1 vccd1 vccd1 _13552_/A sky130_fd_sc_hd__and2_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10763_ _19507_/Q _19121_/Q _19571_/Q _18727_/Q _10650_/S _09482_/A vssd1 vssd1 vccd1
+ vccd1 _10764_/B sky130_fd_sc_hd__mux4_1
XFILLER_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ _12502_/A _12503_/B vssd1 vssd1 vccd1 vccd1 _12502_/Y sky130_fd_sc_hd__nor2_1
X_16270_ _16270_/A vssd1 vssd1 vccd1 vccd1 _16279_/S sky130_fd_sc_hd__buf_6
XFILLER_9_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13482_ _18400_/Q _12598_/B _13486_/S vssd1 vssd1 vccd1 vccd1 _13483_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10694_ _10701_/A _10694_/B vssd1 vssd1 vccd1 vccd1 _10694_/Y sky130_fd_sc_hd__nor2_1
X_15221_ _18676_/Q _15219_/X _15233_/S vssd1 vssd1 vccd1 vccd1 _15222_/A sky130_fd_sc_hd__mux2_1
X_12433_ _19758_/Q _12434_/B vssd1 vssd1 vccd1 vccd1 _12433_/X sky130_fd_sc_hd__or2_1
XANTENNA__11689__A _11776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10593__A _10593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09159__A _11156_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15152_ _16654_/A vssd1 vssd1 vccd1 vccd1 _15152_/X sky130_fd_sc_hd__clkbuf_2
X_12364_ _12294_/S _12362_/Y _12363_/Y _11980_/A vssd1 vssd1 vccd1 vccd1 _12364_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14103_ _14103_/A _14103_/B vssd1 vssd1 vccd1 vccd1 _14103_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__15595__S _15603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17376__A _17376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11315_ _11320_/A _11321_/B _11321_/C vssd1 vssd1 vccd1 vccd1 _11484_/B sky130_fd_sc_hd__and3_1
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15083_ _14553_/A _11619_/Y _15092_/S vssd1 vssd1 vccd1 vccd1 _15083_/X sky130_fd_sc_hd__mux2_1
X_12295_ _19683_/Q _11989_/X _11790_/X vssd1 vssd1 vccd1 vccd1 _12295_/X sky130_fd_sc_hd__o21a_1
XFILLER_141_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14034_ _13760_/X _13770_/X _14034_/S vssd1 vssd1 vccd1 vccd1 _14035_/A sky130_fd_sc_hd__mux2_1
X_18911_ _19337_/CLK _18911_/D vssd1 vssd1 vccd1 vccd1 _18911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11246_ _11242_/B _11083_/Y _11245_/Y vssd1 vssd1 vccd1 vccd1 _11261_/A sky130_fd_sc_hd__a21oi_1
XFILLER_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09752__A1 _09430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18842_ _19590_/CLK _18842_/D vssd1 vssd1 vccd1 vccd1 _18842_/Q sky130_fd_sc_hd__dfxtp_1
X_11177_ _18845_/Q _19399_/Q _19561_/Q _18813_/Q _10185_/S _09736_/A vssd1 vssd1 vccd1
+ vccd1 _11178_/B sky130_fd_sc_hd__mux4_1
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10993__S0 _10909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10128_ _10328_/S vssd1 vssd1 vccd1 vccd1 _10129_/S sky130_fd_sc_hd__buf_4
XFILLER_95_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18773_ _19326_/CLK _18773_/D vssd1 vssd1 vccd1 vccd1 _18773_/Q sky130_fd_sc_hd__dfxtp_1
X_15985_ _16031_/S vssd1 vssd1 vccd1 vccd1 _15994_/S sky130_fd_sc_hd__buf_2
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17315__S _17317_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10059_ _10064_/A _10059_/B vssd1 vssd1 vccd1 vccd1 _10059_/X sky130_fd_sc_hd__or2_1
X_17724_ _17772_/S vssd1 vssd1 vccd1 vccd1 _17724_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14936_ _14838_/X _14935_/X _14898_/X vssd1 vssd1 vccd1 vccd1 _14936_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12967__B _14638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14867_ _16787_/A vssd1 vssd1 vccd1 vccd1 _14867_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17655_ _18468_/Q _17656_/B vssd1 vssd1 vccd1 vccd1 _17667_/C sky130_fd_sc_hd__or2_2
XFILLER_91_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13818_ _13891_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13899_/A sky130_fd_sc_hd__nand2_1
X_16606_ _16606_/A vssd1 vssd1 vccd1 vccd1 _19258_/D sky130_fd_sc_hd__clkbuf_1
X_17586_ _19651_/Q _16816_/A _17590_/S vssd1 vssd1 vccd1 vccd1 _17587_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14798_ _18434_/Q _13228_/B _15051_/S vssd1 vssd1 vccd1 vccd1 _14798_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19325_ _19397_/CLK _19325_/D vssd1 vssd1 vccd1 vccd1 _19325_/Q sky130_fd_sc_hd__dfxtp_1
X_16537_ _16537_/A vssd1 vssd1 vccd1 vccd1 _19225_/D sky130_fd_sc_hd__clkbuf_1
X_13749_ _14034_/S vssd1 vssd1 vccd1 vccd1 _13969_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__12983__A _12983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16455__A _16501_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17050__S _17058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11170__S0 _09692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19256_ _19337_/CLK _19256_/D vssd1 vssd1 vccd1 vccd1 _19256_/Q sky130_fd_sc_hd__dfxtp_1
X_16468_ _16468_/A vssd1 vssd1 vccd1 vccd1 _19194_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13367__A2 _13364_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18207_ _18207_/A _18207_/B vssd1 vssd1 vccd1 vccd1 _19856_/D sky130_fd_sc_hd__nor2_1
X_15419_ _15419_/A vssd1 vssd1 vccd1 vccd1 _18753_/D sky130_fd_sc_hd__clkbuf_1
X_19187_ _19638_/CLK _19187_/D vssd1 vssd1 vccd1 vccd1 _19187_/Q sky130_fd_sc_hd__dfxtp_1
X_16399_ _16399_/A vssd1 vssd1 vccd1 vccd1 _19164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18138_ _18140_/B _18140_/C _18137_/Y vssd1 vssd1 vccd1 vccd1 _19832_/D sky130_fd_sc_hd__o21a_1
XFILLER_117_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10050__A1 _09927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18069_ _18077_/A _18069_/B _18069_/C vssd1 vssd1 vccd1 vccd1 _19809_/D sky130_fd_sc_hd__nor3_1
XANTENNA__10050__B2 _18447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09418__S1 _09364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09911_ _18609_/Q _19298_/Q _09911_/S vssd1 vssd1 vccd1 vccd1 _09911_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09842_ _18611_/Q _19300_/Q _09911_/S vssd1 vssd1 vccd1 vccd1 _09843_/B sky130_fd_sc_hd__mux2_1
XFILLER_113_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _09995_/A vssd1 vssd1 vccd1 vccd1 _10093_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_14_0_clock clkbuf_3_7_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_14_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_39_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11781__B _13630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10678__A _11027_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11161__S0 _09692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17741__A1 _19683_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09207_ _10827_/A vssd1 vssd1 vccd1 vccd1 _09208_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09138_ _10969_/A vssd1 vssd1 vccd1 vccd1 _09139_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_120_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14613__A _14648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11100_ _18830_/Q _19384_/Q _19546_/Q _18798_/Q _10350_/S _09539_/A vssd1 vssd1 vccd1
+ vccd1 _11100_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09707__A _10262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_192_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ _14124_/A _12131_/B _14140_/B vssd1 vssd1 vccd1 vccd1 _12081_/B sky130_fd_sc_hd__nor3_1
XFILLER_104_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14332__B _14332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11031_ _18753_/Q _18982_/Q _18913_/Q _19211_/Q _10959_/X _10960_/X vssd1 vssd1 vccd1
+ vccd1 _11031_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12133__A _14178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15770_ _15770_/A vssd1 vssd1 vccd1 vccd1 _18895_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _18308_/Q _12982_/B _12982_/C vssd1 vssd1 vccd1 vccd1 _12983_/C sky130_fd_sc_hd__and3_1
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13294__B2 _18633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10727__S0 _10724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _15010_/A vssd1 vssd1 vccd1 vccd1 _15077_/S sky130_fd_sc_hd__buf_8
XANTENNA_input12_A io_dbus_rdata[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09442__A _09538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ _12119_/S _11957_/B _11932_/X _14431_/B vssd1 vssd1 vccd1 vccd1 _11933_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_91_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _16813_/X _19586_/Q _17446_/S vssd1 vssd1 vccd1 vccd1 _17441_/A sky130_fd_sc_hd__mux2_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _14652_/A vssd1 vssd1 vccd1 vccd1 _18570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11864_ _11939_/A vssd1 vssd1 vccd1 vccd1 _14005_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _13603_/A vssd1 vssd1 vccd1 vccd1 _14138_/B sky130_fd_sc_hd__buf_2
XFILLER_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17371_ _17371_/A vssd1 vssd1 vccd1 vccd1 _19555_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _09169_/A _10814_/X _09177_/A vssd1 vssd1 vccd1 vccd1 _10815_/X sky130_fd_sc_hd__a21o_1
X_14583_ _11517_/B _14526_/B _14582_/Y _14573_/X vssd1 vssd1 vccd1 vccd1 _18550_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11795_ _11787_/Y _11794_/Y _12165_/S vssd1 vssd1 vccd1 vccd1 _11795_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19110_ _19723_/CLK _19110_/D vssd1 vssd1 vccd1 vccd1 _19110_/Q sky130_fd_sc_hd__dfxtp_1
X_16322_ _16322_/A vssd1 vssd1 vccd1 vccd1 _19130_/D sky130_fd_sc_hd__clkbuf_1
X_13534_ _13542_/A _13534_/B vssd1 vssd1 vccd1 vccd1 _13535_/A sky130_fd_sc_hd__and2_1
XFILLER_159_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10746_ _19409_/Q _19185_/Q _19702_/Q _19153_/Q _10858_/A _10740_/X vssd1 vssd1 vccd1
+ vccd1 _10746_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17732__A1 _19681_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19041_ _19723_/CLK _19041_/D vssd1 vssd1 vccd1 vccd1 _19041_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13411__B _13411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16253_ _16090_/X _19100_/Q _16257_/S vssd1 vssd1 vccd1 vccd1 _16254_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13465_ _13465_/A vssd1 vssd1 vccd1 vccd1 _18392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10677_ _10983_/S vssd1 vssd1 vccd1 vccd1 _11027_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__12308__A _14265_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15204_ _15220_/A vssd1 vssd1 vccd1 vccd1 _15217_/S sky130_fd_sc_hd__buf_4
XFILLER_145_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12416_ _12439_/B _12415_/Y _11859_/X vssd1 vssd1 vccd1 vccd1 _12416_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16184_ _16184_/A vssd1 vssd1 vccd1 vccd1 _19065_/D sky130_fd_sc_hd__clkbuf_1
X_13396_ _13067_/B _13178_/X _12665_/A _18102_/B _13395_/X vssd1 vssd1 vccd1 vccd1
+ _13396_/X sky130_fd_sc_hd__a221o_1
XFILLER_127_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09973__A1 _09927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15135_ _16430_/A _16357_/B _15412_/C vssd1 vssd1 vccd1 vccd1 _17463_/A sky130_fd_sc_hd__or3_4
XANTENNA__09973__B2 _18448_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12347_ _12419_/A _12347_/B vssd1 vssd1 vccd1 vccd1 _14289_/A sky130_fd_sc_hd__nand2_4
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output80_A _12096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15066_ _16841_/A vssd1 vssd1 vccd1 vccd1 _15066_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12278_ _12277_/Y _12173_/Y _11831_/X _12497_/A vssd1 vssd1 vccd1 vccd1 _12280_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_14017_ _13692_/X _13629_/X _14034_/S vssd1 vssd1 vccd1 vccd1 _14018_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11229_ _11229_/A vssd1 vssd1 vccd1 vccd1 _11229_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12043__A _12043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11532__A1 _14543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__S0 _10664_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18825_ _19539_/CLK _18825_/D vssd1 vssd1 vccd1 vccd1 _18825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17045__S _17047_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11882__A _11901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18756_ _19597_/CLK _18756_/D vssd1 vssd1 vccd1 vccd1 _18756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15968_ _14740_/X _18984_/Q _15972_/S vssd1 vssd1 vccd1 vccd1 _15969_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09352__A _09352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17707_ _17707_/A vssd1 vssd1 vccd1 vccd1 _17708_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14919_ _14918_/X _18603_/Q _14941_/S vssd1 vssd1 vccd1 vccd1 _14920_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18687_ _19779_/CLK _18687_/D vssd1 vssd1 vccd1 vccd1 _18687_/Q sky130_fd_sc_hd__dfxtp_1
X_15899_ _15899_/A vssd1 vssd1 vccd1 vccd1 _18952_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17638_ _17638_/A vssd1 vssd1 vccd1 vccd1 _19665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17569_ _17569_/A vssd1 vssd1 vccd1 vccd1 _19643_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09887__S1 _09881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19308_ _19691_/CLK _19308_/D vssd1 vssd1 vccd1 vccd1 _19308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19239_ _19625_/CLK _19239_/D vssd1 vssd1 vccd1 vccd1 _19239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09639__S1 _09695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12012__A2 _14093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15529__A _16784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14433__A _14591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11771__A1 _17762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09527__A _10496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09811__S1 _09810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10957__S0 _10909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _18610_/Q _19299_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09826_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input4_A io_dbus_rdata[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11792__A _19733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09756_ _09756_/A _09756_/B _11224_/A vssd1 vssd1 vccd1 vccd1 _11152_/C sky130_fd_sc_hd__and3_1
XFILLER_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09687_ _09688_/A _12501_/A vssd1 vssd1 vccd1 vccd1 _09901_/A sky130_fd_sc_hd__and2_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17411__A0 _16771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15017__A2 _14958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_139_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11016__B _11016_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10600_ _10601_/B _12474_/B vssd1 vssd1 vccd1 vccd1 _11244_/A sky130_fd_sc_hd__and2b_1
XFILLER_120_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11580_ _11736_/A _11592_/A _11580_/C _11599_/B vssd1 vssd1 vccd1 vccd1 _11580_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10531_ _19639_/Q _19056_/Q _19093_/Q _18699_/Q _10560_/S _09634_/A vssd1 vssd1 vccd1
+ vccd1 _10531_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13250_ _19479_/Q _13235_/X _13236_/X _18360_/Q _13249_/X vssd1 vssd1 vccd1 vccd1
+ _13253_/A sky130_fd_sc_hd__a221o_1
XFILLER_109_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10462_ _10462_/A _10462_/B vssd1 vssd1 vccd1 vccd1 _11242_/A sky130_fd_sc_hd__and2_1
XFILLER_109_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12201_ _19748_/Q _12186_/X _12194_/X _12200_/X vssd1 vssd1 vccd1 vccd1 _12201_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_129_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15439__A _15485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13181_ _18623_/Q _13181_/B vssd1 vssd1 vccd1 vccd1 _13181_/X sky130_fd_sc_hd__or2_1
XFILLER_124_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10393_ _18767_/Q _18996_/Q _18927_/Q _19225_/Q _10230_/X _11111_/A vssd1 vssd1 vccd1
+ vccd1 _10394_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09437__A _10982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ _12348_/A _12132_/B vssd1 vssd1 vccd1 vccd1 _12133_/B sky130_fd_sc_hd__nand2_1
XFILLER_150_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16969__S _16975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16940_ _16771_/X _19379_/Q _16942_/S vssd1 vssd1 vccd1 vccd1 _16941_/A sky130_fd_sc_hd__mux2_1
X_12063_ _12063_/A _13603_/A vssd1 vssd1 vccd1 vccd1 _12064_/B sky130_fd_sc_hd__nor2_1
XFILLER_104_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11014_ _11060_/A _11014_/B vssd1 vssd1 vccd1 vccd1 _11014_/X sky130_fd_sc_hd__or2_1
X_16871_ _16917_/S vssd1 vssd1 vccd1 vccd1 _16880_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18610_ _19395_/CLK _18610_/D vssd1 vssd1 vccd1 vccd1 _18610_/Q sky130_fd_sc_hd__dfxtp_1
X_15822_ _14772_/X _18918_/Q _15830_/S vssd1 vssd1 vccd1 vccd1 _15823_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19590_ _19590_/CLK _19590_/D vssd1 vssd1 vccd1 vccd1 _19590_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09172__A _09172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18541_ _18548_/CLK _18541_/D vssd1 vssd1 vccd1 vccd1 _18541_/Q sky130_fd_sc_hd__dfxtp_1
X_15753_ _15753_/A vssd1 vssd1 vccd1 vccd1 _18887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ _18225_/A vssd1 vssd1 vccd1 vccd1 _14673_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17402__A0 _16758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10176__S1 _09723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11916_ _10554_/B _18500_/Q _11948_/A vssd1 vssd1 vccd1 vccd1 _13622_/A sky130_fd_sc_hd__mux2_2
X_14704_ _19081_/Q vssd1 vssd1 vccd1 vccd1 _14922_/S sky130_fd_sc_hd__buf_2
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15684_ _18857_/Q _15516_/X _15686_/S vssd1 vssd1 vccd1 vccd1 _15685_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18472_ _19080_/CLK _18472_/D vssd1 vssd1 vccd1 vccd1 _18472_/Q sky130_fd_sc_hd__dfxtp_1
X_12896_ _12933_/C vssd1 vssd1 vccd1 vccd1 _12897_/B sky130_fd_sc_hd__buf_2
XFILLER_166_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _14654_/A _14635_/B vssd1 vssd1 vccd1 vccd1 _14636_/A sky130_fd_sc_hd__and2_1
XFILLER_33_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15964__A0 _14714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17423_ _17423_/A vssd1 vssd1 vccd1 vccd1 _19578_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _14431_/B vssd1 vssd1 vccd1 vccd1 _11847_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16209__S _16209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13422__A _18649_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _17376_/A vssd1 vssd1 vccd1 vccd1 _17363_/S sky130_fd_sc_hd__buf_4
X_14566_ _14566_/A _14580_/B vssd1 vssd1 vccd1 vccd1 _14566_/X sky130_fd_sc_hd__or2_1
XFILLER_60_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11778_ _13939_/B _11778_/B vssd1 vssd1 vccd1 vccd1 _11811_/A sky130_fd_sc_hd__xnor2_1
X_16305_ _16061_/X _19123_/Q _16307_/S vssd1 vssd1 vccd1 vccd1 _16306_/A sky130_fd_sc_hd__mux2_1
X_13517_ _13563_/A vssd1 vssd1 vccd1 vccd1 _13542_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17829__A _17840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10729_ _10803_/A _10727_/X _10728_/X vssd1 vssd1 vccd1 vccd1 _10729_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10257__S _10257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17285_ _19517_/Q _16693_/X _17291_/S vssd1 vssd1 vccd1 vccd1 _17286_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14497_ _14497_/A vssd1 vssd1 vccd1 vccd1 _18518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19024_ _19444_/CLK _19024_/D vssd1 vssd1 vccd1 vccd1 _19024_/Q sky130_fd_sc_hd__dfxtp_1
X_16236_ _16236_/A vssd1 vssd1 vccd1 vccd1 _19092_/D sky130_fd_sc_hd__clkbuf_1
X_13448_ _13448_/A vssd1 vssd1 vccd1 vccd1 _18384_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15192__A1 _15191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16167_ _16167_/A vssd1 vssd1 vccd1 vccd1 _19057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13379_ _13390_/A _18646_/Q vssd1 vssd1 vccd1 vccd1 _13379_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11753__A1 _19731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15118_ _15125_/A vssd1 vssd1 vccd1 vccd1 _15118_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11596__B _12510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16098_ _16098_/A vssd1 vssd1 vccd1 vccd1 _19033_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11088__S _11088_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15783__S _15791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15049_ _18487_/Q _15049_/B vssd1 vssd1 vccd1 vccd1 _15059_/B sky130_fd_sc_hd__and2_1
XFILLER_141_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19857_ _19858_/CLK _19857_/D vssd1 vssd1 vccd1 vccd1 _19857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09610_ _09610_/A vssd1 vssd1 vccd1 vccd1 _09610_/X sky130_fd_sc_hd__clkbuf_4
X_18808_ _19556_/CLK _18808_/D vssd1 vssd1 vccd1 vccd1 _18808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19788_ _19788_/CLK _19788_/D vssd1 vssd1 vccd1 vccd1 _19788_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12501__A _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09541_ _10306_/A vssd1 vssd1 vccd1 vccd1 _09542_/A sky130_fd_sc_hd__buf_2
X_18739_ _19714_/CLK _18739_/D vssd1 vssd1 vccd1 vccd1 _18739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17503__S _17507_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09472_ _10844_/A vssd1 vssd1 vccd1 vccd1 _10895_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_140_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09810__A _09810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10956__A _10956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15023__S _15056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10244__A1 _10239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19579_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13478__S _13486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14163__A _14163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_65_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13497__A1 _12779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10704__C1 _10944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09808_ _09808_/A vssd1 vssd1 vccd1 vccd1 _09872_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_47_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09739_ _11178_/A _09738_/X _09317_/A vssd1 vssd1 vccd1 vccd1 _09739_/X sky130_fd_sc_hd__o21a_1
XANTENNA__18188__A1 _19850_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12130__B _14168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10158__S1 _09145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17413__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12750_ _12830_/B _12525_/X _12749_/X _19815_/Q vssd1 vssd1 vccd1 vccd1 _12750_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11652_/X _11655_/B _11653_/A vssd1 vssd1 vccd1 vccd1 _11702_/B sky130_fd_sc_hd__a21o_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12681_ _19795_/Q _12665_/X _12666_/X _12679_/X _12680_/X vssd1 vssd1 vccd1 vccd1
+ _12681_/X sky130_fd_sc_hd__a221o_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10483__B2 _18437_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16029__S _16031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14420_/A vssd1 vssd1 vccd1 vccd1 _18485_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11688_/C vssd1 vssd1 vccd1 vccd1 _13789_/A sky130_fd_sc_hd__inv_2
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14057__B _14057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17699__A0 _19676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15868__S _15874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14351_ _18462_/Q vssd1 vssd1 vccd1 vccd1 _14765_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11563_ _12412_/B vssd1 vssd1 vccd1 vccd1 _11563_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13302_ _18282_/Q _13126_/X _13127_/X _18365_/Q vssd1 vssd1 vccd1 vccd1 _13302_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17070_ _17070_/A vssd1 vssd1 vccd1 vccd1 _19436_/D sky130_fd_sc_hd__clkbuf_1
X_10514_ _19413_/Q _19189_/Q _19706_/Q _19157_/Q _10500_/X _10501_/X vssd1 vssd1 vccd1
+ vccd1 _10514_/X sky130_fd_sc_hd__mux4_1
X_14282_ _18452_/Q _14281_/X _14306_/S vssd1 vssd1 vccd1 vccd1 _14283_/A sky130_fd_sc_hd__mux2_1
X_11494_ _18561_/Q vssd1 vssd1 vccd1 vccd1 _11511_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_171_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16021_ _15022_/X _19008_/Q _16027_/S vssd1 vssd1 vccd1 vccd1 _16022_/A sky130_fd_sc_hd__mux2_1
X_13233_ _13185_/X _13230_/X _13231_/X _13232_/X vssd1 vssd1 vccd1 vccd1 _18358_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10445_ _10219_/X _10438_/Y _10440_/Y _10442_/Y _10444_/Y vssd1 vssd1 vccd1 vccd1
+ _10445_/X sky130_fd_sc_hd__o32a_1
XFILLER_136_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11735__A1 _14559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13164_ _12556_/X _13152_/Y _13163_/X _12712_/X _18621_/Q vssd1 vssd1 vccd1 vccd1
+ _15254_/B sky130_fd_sc_hd__a32oi_4
XFILLER_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10376_ _19643_/Q _19060_/Q _19097_/Q _18703_/Q _09448_/S _09554_/A vssd1 vssd1 vccd1
+ vccd1 _10376_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12115_ _14163_/A vssd1 vssd1 vccd1 vccd1 _12115_/Y sky130_fd_sc_hd__inv_2
X_17972_ _17980_/A _17972_/B _17973_/B vssd1 vssd1 vccd1 vccd1 _19775_/D sky130_fd_sc_hd__nor3_1
X_13095_ _14601_/A vssd1 vssd1 vccd1 vccd1 _17892_/A sky130_fd_sc_hd__buf_4
XANTENNA__14801__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19711_ _19714_/CLK _19711_/D vssd1 vssd1 vccd1 vccd1 _19711_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09787__S0 _09760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12046_ _12072_/A vssd1 vssd1 vccd1 vccd1 _17204_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16923_ _16743_/X _19371_/Q _16931_/S vssd1 vssd1 vccd1 vccd1 _16924_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19642_ _19642_/CLK _19642_/D vssd1 vssd1 vccd1 vccd1 _19642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16854_ _19341_/Q _16648_/X _16858_/S vssd1 vssd1 vccd1 vccd1 _16855_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _15805_/A vssd1 vssd1 vccd1 vccd1 _18911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19573_ _19704_/CLK _19573_/D vssd1 vssd1 vccd1 vccd1 _19573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13997_ _13888_/X _13884_/X _13997_/S vssd1 vssd1 vccd1 vccd1 _14135_/B sky130_fd_sc_hd__mux2_1
X_16785_ _16784_/X _19319_/Q _16791_/S vssd1 vssd1 vccd1 vccd1 _16786_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16728__A _16728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18524_ _19733_/CLK _18524_/D vssd1 vssd1 vccd1 vccd1 _18524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12948_ _17895_/A vssd1 vssd1 vccd1 vccd1 _12948_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15736_ _17391_/A _17463_/A vssd1 vssd1 vccd1 vccd1 _15793_/A sky130_fd_sc_hd__or2_2
XFILLER_34_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18455_ _19081_/CLK _18455_/D vssd1 vssd1 vccd1 vccd1 _18455_/Q sky130_fd_sc_hd__dfxtp_4
X_12879_ _18273_/Q vssd1 vssd1 vccd1 vccd1 _12883_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15667_ _18849_/Q _15487_/X _15675_/S vssd1 vssd1 vccd1 vccd1 _15668_/A sky130_fd_sc_hd__mux2_1
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17406_ _17406_/A vssd1 vssd1 vccd1 vccd1 _19570_/D sky130_fd_sc_hd__clkbuf_1
X_14618_ _14638_/A _14618_/B vssd1 vssd1 vccd1 vccd1 _18560_/D sky130_fd_sc_hd__nor2_1
X_18386_ _18386_/CLK _18386_/D vssd1 vssd1 vccd1 vccd1 _18386_/Q sky130_fd_sc_hd__dfxtp_1
X_15598_ _15598_/A vssd1 vssd1 vccd1 vccd1 _18818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15778__S _15780_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09711__S0 _10257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14549_ _18536_/Q _14522_/X _14547_/Y _14548_/X vssd1 vssd1 vccd1 vccd1 _18536_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17337_ _16768_/X _19540_/Q _17341_/S vssd1 vssd1 vccd1 vccd1 _17338_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17559__A _17605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12991__A _12991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11974__A1 _18502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17268_ _17268_/A vssd1 vssd1 vccd1 vccd1 _19509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19007_ _19331_/CLK _19007_/D vssd1 vssd1 vccd1 vccd1 _19007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16219_ _16219_/A vssd1 vssd1 vccd1 vccd1 _19084_/D sky130_fd_sc_hd__clkbuf_1
X_17199_ _19486_/Q _17198_/X _17206_/S vssd1 vssd1 vccd1 vccd1 _17200_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12923__B1 _12922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12215__B _19748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16402__S _16402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14711__A _14842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10450__S _10450_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09524_ _10395_/A _09524_/B vssd1 vssd1 vccd1 vccd1 _09524_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16357__B _16357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09540__A _09554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_141_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _18509_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _19433_/Q _19209_/Q _19726_/Q _19177_/Q _10465_/S _09442_/X vssd1 vssd1 vccd1
+ vccd1 _09455_/X sky130_fd_sc_hd__mux4_1
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09386_ _19434_/Q _19210_/Q _19727_/Q _19178_/Q _09369_/S _09364_/A vssd1 vssd1 vccd1
+ vccd1 _09386_/X sky130_fd_sc_hd__mux4_2
XANTENNA__09607__B1 _09394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11965__A1 _19739_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_156_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19698_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10312__S1 _09555_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11717__A1 _11822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10230_ _10486_/S vssd1 vssd1 vccd1 vccd1 _10230_/X sky130_fd_sc_hd__buf_4
XFILLER_145_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10161_ _10007_/A _10152_/X _10156_/X _10160_/X _09135_/A vssd1 vssd1 vccd1 vccd1
+ _10161_/X sky130_fd_sc_hd__a311o_1
XFILLER_161_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16312__S _16318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10555__A_N _10554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10092_ _18837_/Q _19391_/Q _19553_/Q _18805_/Q _10153_/S _09769_/A vssd1 vssd1 vccd1
+ vccd1 _10093_/B sky130_fd_sc_hd__mux4_1
XFILLER_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11456__S _14120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13920_ _13918_/S _13919_/X _13819_/X vssd1 vssd1 vccd1 vccd1 _14293_/B sky130_fd_sc_hd__o21ai_1
XFILLER_59_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13851_ _13837_/X _13842_/Y _13850_/X _13810_/A vssd1 vssd1 vccd1 vccd1 _13851_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15092__A0 _14559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12802_ _18173_/A vssd1 vssd1 vccd1 vccd1 _12802_/X sky130_fd_sc_hd__buf_4
XANTENNA__17143__S _17143_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13782_ _13752_/X _13763_/X _13780_/X _14122_/S vssd1 vssd1 vccd1 vccd1 _13782_/X
+ sky130_fd_sc_hd__o22a_1
X_16570_ _16570_/A vssd1 vssd1 vccd1 vccd1 _19240_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13642__A1 _12424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10994_ _10956_/A _10993_/X _10827_/A vssd1 vssd1 vccd1 vccd1 _10994_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_109_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _18381_/CLK sky130_fd_sc_hd__clkbuf_16
X_12733_ _13426_/A _18642_/Q vssd1 vssd1 vccd1 vccd1 _12733_/Y sky130_fd_sc_hd__nand2_1
X_15521_ _15521_/A vssd1 vssd1 vccd1 vccd1 _18794_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09941__S0 _09866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16982__S _16986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18240_ _18239_/B _18239_/C _19868_/Q vssd1 vssd1 vccd1 vccd1 _18241_/C sky130_fd_sc_hd__a21oi_1
XFILLER_30_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15452_ _15452_/A vssd1 vssd1 vccd1 vccd1 _18768_/D sky130_fd_sc_hd__clkbuf_1
X_12664_ _12664_/A vssd1 vssd1 vccd1 vccd1 _12665_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _18480_/Q vssd1 vssd1 vccd1 vccd1 _17728_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11615_ _12460_/A _11831_/A _11614_/X vssd1 vssd1 vccd1 vccd1 _11688_/C sky130_fd_sc_hd__a21oi_4
X_18171_ _19844_/Q _18175_/C _18170_/X vssd1 vssd1 vccd1 vccd1 _18171_/Y sky130_fd_sc_hd__a21oi_1
X_15383_ _15383_/A vssd1 vssd1 vccd1 vccd1 _18739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12595_ _12712_/A vssd1 vssd1 vccd1 vccd1 _13306_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17122_ _16825_/X _19460_/Q _17130_/S vssd1 vssd1 vccd1 vccd1 _17123_/A sky130_fd_sc_hd__mux2_1
X_14334_ _14331_/A _13975_/X _13721_/X _14333_/X vssd1 vssd1 vccd1 vccd1 _14334_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__13700__A _13711_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11546_ _19081_/Q vssd1 vssd1 vccd1 vccd1 _15060_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17053_ _17053_/A vssd1 vssd1 vccd1 vccd1 _19429_/D sky130_fd_sc_hd__clkbuf_1
X_14265_ _14265_/A _14265_/B vssd1 vssd1 vccd1 vccd1 _14265_/Y sky130_fd_sc_hd__nor2_1
XFILLER_167_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11477_ _11477_/A _11587_/A vssd1 vssd1 vccd1 vccd1 _11482_/B sky130_fd_sc_hd__nor2_1
XFILLER_171_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16004_ _16004_/A vssd1 vssd1 vccd1 vccd1 _19000_/D sky130_fd_sc_hd__clkbuf_1
X_13216_ _13110_/A _13118_/X _13215_/X _13167_/X vssd1 vssd1 vccd1 vccd1 _18357_/D
+ sky130_fd_sc_hd__o211a_1
X_10428_ _10428_/A _10428_/B vssd1 vssd1 vccd1 vccd1 _10428_/X sky130_fd_sc_hd__or2_1
X_14196_ _13594_/X _14087_/X _14195_/X _14097_/X vssd1 vssd1 vccd1 vccd1 _14196_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10916__C1 _09223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12035__B _13607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13147_ _19761_/Q _13123_/A _13143_/X _13146_/X vssd1 vssd1 vccd1 vccd1 _13148_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_125_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16222__S _16224_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10359_ _10752_/A vssd1 vssd1 vccd1 vccd1 _10566_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14531__A _15134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09625__A _09625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17955_ _17980_/A _17955_/B _17955_/C vssd1 vssd1 vccd1 vccd1 _19769_/D sky130_fd_sc_hd__nor3_1
X_13078_ _18348_/Q _15242_/A vssd1 vssd1 vccd1 vccd1 _13078_/X sky130_fd_sc_hd__and2_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16906_ _16906_/A vssd1 vssd1 vccd1 vccd1 _19364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12029_ _12131_/A vssd1 vssd1 vccd1 vccd1 _14124_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12051__A _13295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17886_ _17886_/A vssd1 vssd1 vccd1 vccd1 _17886_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12684__A2 _18622_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19625_ _19625_/CLK _19625_/D vssd1 vssd1 vccd1 vccd1 _19625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16837_ _16837_/A vssd1 vssd1 vccd1 vccd1 _19335_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12986__A _12997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15083__A0 _14553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19556_ _19556_/CLK _19556_/D vssd1 vssd1 vccd1 vccd1 _19556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12436__A2 _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13633__A1 _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16768_ _16768_/A vssd1 vssd1 vccd1 vccd1 _16768_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09360__A _10132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18507_ _18510_/CLK _18507_/D vssd1 vssd1 vccd1 vccd1 _18507_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09932__S0 _09874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15719_ _18873_/Q _15567_/X _15719_/S vssd1 vssd1 vccd1 vccd1 _15720_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19487_ _19488_/CLK _19487_/D vssd1 vssd1 vccd1 vccd1 _19487_/Q sky130_fd_sc_hd__dfxtp_1
X_16699_ _16699_/A vssd1 vssd1 vccd1 vccd1 _16699_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09240_ _09856_/A _09240_/B vssd1 vssd1 vccd1 vccd1 _09240_/X sky130_fd_sc_hd__or2_1
X_18438_ _19078_/CLK _18438_/D vssd1 vssd1 vccd1 vccd1 _18438_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_167_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_73_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19716_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_147_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09171_ _09171_/A vssd1 vssd1 vccd1 vccd1 _09172_/A sky130_fd_sc_hd__clkbuf_4
X_18369_ _18402_/CLK _18369_/D vssd1 vssd1 vccd1 vccd1 _18369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_88_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19795_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__16921__A _16977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14897__A0 _18442_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11130__A _11130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09999__S0 _09976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16132__S _16135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_11_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19592_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09535__A _09640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10979__A2_N _11070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11883__A0 _11880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_26_clock clkbuf_opt_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19647_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13624__A1 _13623_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09507_ _10762_/A vssd1 vssd1 vccd1 vccd1 _10638_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _10733_/S vssd1 vssd1 vccd1 vccd1 _09629_/A sky130_fd_sc_hd__clkbuf_4
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11024__B _12460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09369_ _18617_/Q _19306_/Q _09369_/S vssd1 vssd1 vccd1 vccd1 _09370_/B sky130_fd_sc_hd__mux2_1
XFILLER_138_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11938__A1 _11984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15211__S _15217_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11400_ _11400_/A vssd1 vssd1 vccd1 vccd1 _12520_/A sky130_fd_sc_hd__buf_2
XFILLER_165_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15129__B2 _11199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12380_ _11199_/A _18518_/Q _12423_/S vssd1 vssd1 vccd1 vccd1 _12381_/A sky130_fd_sc_hd__mux2_8
XFILLER_165_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10071__C1 _09395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ _18580_/Q _18579_/Q vssd1 vssd1 vccd1 vccd1 _11519_/B sky130_fd_sc_hd__or2_2
XANTENNA__17927__A _19761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14050_ _11899_/Y _13730_/X _14049_/X vssd1 vssd1 vccd1 vccd1 _14050_/X sky130_fd_sc_hd__a21bo_1
X_11262_ _11262_/A _11262_/B vssd1 vssd1 vccd1 vccd1 _11263_/B sky130_fd_sc_hd__nor2_1
X_13001_ _13003_/B _13003_/C _13000_/Y vssd1 vssd1 vccd1 vccd1 _18313_/D sky130_fd_sc_hd__o21a_1
X_10213_ _18834_/Q _19388_/Q _19550_/Q _18802_/Q _09795_/A _10080_/X vssd1 vssd1 vccd1
+ vccd1 _10213_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11193_ _10327_/A _11192_/X _09621_/A vssd1 vssd1 vccd1 vccd1 _11193_/X sky130_fd_sc_hd__o21a_1
XFILLER_161_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input42_A io_ibus_inst[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09445__A _09629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10144_ _10144_/A _10144_/B vssd1 vssd1 vccd1 vccd1 _10144_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17740_ _17730_/X _12779_/X _17724_/X vssd1 vssd1 vccd1 vccd1 _17740_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10075_ _18606_/Q _19295_/Q _10075_/S vssd1 vssd1 vccd1 vccd1 _10075_/X sky130_fd_sc_hd__mux2_1
X_14952_ _15010_/A vssd1 vssd1 vccd1 vccd1 _14997_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_75_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13903_ _14212_/A _13667_/X _13797_/X _13902_/X vssd1 vssd1 vccd1 vccd1 _13903_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10221__S0 _09673_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17671_ _19671_/Q _17670_/X _17681_/S vssd1 vssd1 vccd1 vccd1 _17672_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14883_ _14883_/A _14894_/C vssd1 vssd1 vccd1 vccd1 _14883_/Y sky130_fd_sc_hd__nand2_1
X_19410_ _19506_/CLK _19410_/D vssd1 vssd1 vccd1 vccd1 _19410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16622_ _16622_/A vssd1 vssd1 vccd1 vccd1 _19266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13834_ _13743_/S _13683_/X _13833_/X vssd1 vssd1 vccd1 vccd1 _13964_/A sky130_fd_sc_hd__o21ai_2
XFILLER_90_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19341_ _19633_/CLK _19341_/D vssd1 vssd1 vccd1 vccd1 _19341_/Q sky130_fd_sc_hd__dfxtp_1
X_16553_ _16553_/A vssd1 vssd1 vccd1 vccd1 _19232_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13765_ _13609_/X _13597_/X _13765_/S vssd1 vssd1 vccd1 vccd1 _13765_/X sky130_fd_sc_hd__mux2_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10977_ _10823_/A _10965_/X _10971_/Y _10976_/X vssd1 vssd1 vccd1 vccd1 _10977_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_187_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17601__S _17601_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15504_ _18789_/Q _15503_/X _15504_/S vssd1 vssd1 vccd1 vccd1 _15505_/A sky130_fd_sc_hd__mux2_1
X_12716_ _13106_/B _12713_/X _12714_/X _13516_/B _18299_/Q vssd1 vssd1 vccd1 vccd1
+ _12716_/X sky130_fd_sc_hd__o32a_1
X_19272_ _19559_/CLK _19272_/D vssd1 vssd1 vccd1 vccd1 _19272_/Q sky130_fd_sc_hd__dfxtp_1
X_16484_ _16109_/X _19202_/Q _16486_/S vssd1 vssd1 vccd1 vccd1 _16485_/A sky130_fd_sc_hd__mux2_1
X_13696_ _13656_/X _13693_/X _14086_/S vssd1 vssd1 vccd1 vccd1 _13696_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18223_ _18223_/A _18223_/B vssd1 vssd1 vccd1 vccd1 _18223_/Y sky130_fd_sc_hd__nor2_1
X_12647_ _18336_/Q _12568_/X _13127_/A _13322_/A _12646_/X vssd1 vssd1 vccd1 vccd1
+ _12647_/X sky130_fd_sc_hd__a221o_1
X_15435_ _18761_/Q _15165_/X _15437_/S vssd1 vssd1 vccd1 vccd1 _15436_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18154_ _19838_/Q _18156_/C _18153_/Y vssd1 vssd1 vccd1 vccd1 _19838_/D sky130_fd_sc_hd__o21a_1
XFILLER_156_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15366_ _15366_/A vssd1 vssd1 vccd1 vccd1 _18731_/D sky130_fd_sc_hd__clkbuf_1
X_12578_ _12766_/A vssd1 vssd1 vccd1 vccd1 _13415_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11869__B _13617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10062__C1 _09404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17105_ _17105_/A vssd1 vssd1 vccd1 vccd1 _19452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14317_ _12408_/B _13933_/A _14316_/X _14120_/A vssd1 vssd1 vccd1 vccd1 _14317_/X
+ sky130_fd_sc_hd__o211a_4
X_11529_ _12505_/B _13527_/B _13529_/A _11599_/B vssd1 vssd1 vccd1 vccd1 _11530_/C
+ sky130_fd_sc_hd__and4_1
X_18085_ _18085_/A vssd1 vssd1 vccd1 vccd1 _18120_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15297_ _15297_/A vssd1 vssd1 vccd1 vccd1 _18701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17036_ _19422_/Q _16702_/X _17036_/S vssd1 vssd1 vccd1 vccd1 _17037_/A sky130_fd_sc_hd__mux2_1
X_14248_ _14248_/A vssd1 vssd1 vccd1 vccd1 _18449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14179_ _13796_/A _14180_/B _14177_/X _14178_/X vssd1 vssd1 vccd1 vccd1 _14179_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14261__A _14265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09355__A _10384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18987_ _19569_/CLK _18987_/D vssd1 vssd1 vccd1 vccd1 _18987_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16887__S _16891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15791__S _15791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _17948_/A _17944_/C vssd1 vssd1 vccd1 vccd1 _17938_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10117__B1 _09996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17045__A1 _16715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17869_ _17869_/A vssd1 vssd1 vccd1 vccd1 _19735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13605__A _13643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19608_ _19608_/CLK _19608_/D vssd1 vssd1 vccd1 vccd1 _19608_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10763__S1 _09482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13606__A1 _14155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19539_ _19539_/CLK _19539_/D vssd1 vssd1 vccd1 vccd1 _19539_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09286__B2 _18457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09223_ _09223_/A vssd1 vssd1 vccd1 vccd1 _09224_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14031__A1 _11880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09154_ _10604_/S vssd1 vssd1 vccd1 vccd1 _10466_/S sky130_fd_sc_hd__buf_2
XFILLER_147_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14155__B _14155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_10_0_clock clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_10_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__15966__S _15972_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ _11320_/A _18558_/Q _11321_/B vssd1 vssd1 vccd1 vccd1 _12471_/B sky130_fd_sc_hd__or3b_4
XFILLER_147_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13486__S _13486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09987_ _19425_/Q _19201_/Q _19718_/Q _19169_/Q _09983_/X _09984_/X vssd1 vssd1 vccd1
+ vccd1 _09987_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10659__B2 _10658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10754__S1 _10740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ _19599_/Q _19437_/Q _18883_/Q _18653_/Q _10724_/X _10713_/X vssd1 vssd1 vccd1
+ vccd1 _10900_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11880_ _11880_/A vssd1 vssd1 vccd1 vccd1 _11880_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10831_ _19601_/Q _19439_/Q _18885_/Q _18655_/Q _09152_/A _10740_/A vssd1 vssd1 vccd1
+ vccd1 _10831_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13234__B _18628_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14270__A1 _12313_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13550_ _09106_/Y _13536_/X _13537_/X _14900_/A vssd1 vssd1 vccd1 vccd1 _13551_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12281__A0 _11148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10762_ _10762_/A _10762_/B vssd1 vssd1 vccd1 vccd1 _10762_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12501_ _12501_/A _12503_/B vssd1 vssd1 vccd1 vccd1 _12501_/Y sky130_fd_sc_hd__nor2_1
XFILLER_157_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13481_ _13481_/A vssd1 vssd1 vccd1 vccd1 _18399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16037__S _16049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10693_ _19508_/Q _19122_/Q _19572_/Q _18728_/Q _10770_/S _09512_/A vssd1 vssd1 vccd1
+ vccd1 _10694_/B sky130_fd_sc_hd__mux4_1
XFILLER_13_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12033__A0 _10412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15220_ _15220_/A vssd1 vssd1 vccd1 vccd1 _15233_/S sky130_fd_sc_hd__clkbuf_8
X_12432_ _14319_/A vssd1 vssd1 vccd1 vccd1 _12432_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11689__B _13996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15151_ _15151_/A vssd1 vssd1 vccd1 vccd1 _18654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15876__S _15878_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12363_ _12452_/S _14284_/A vssd1 vssd1 vccd1 vccd1 _12363_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14102_ _14102_/A vssd1 vssd1 vccd1 vccd1 _14102_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09874__S _09874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11314_ _11314_/A _11599_/A vssd1 vssd1 vccd1 vccd1 _11736_/B sky130_fd_sc_hd__or2b_1
X_15082_ _15082_/A vssd1 vssd1 vccd1 vccd1 _18619_/D sky130_fd_sc_hd__clkbuf_1
X_12294_ _12290_/X _12293_/Y _12294_/S vssd1 vssd1 vccd1 vccd1 _12294_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14033_ _14033_/A vssd1 vssd1 vccd1 vccd1 _18434_/D sky130_fd_sc_hd__clkbuf_1
X_18910_ _19725_/CLK _18910_/D vssd1 vssd1 vccd1 vccd1 _18910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11245_ _10557_/A _11247_/B _11081_/A vssd1 vssd1 vccd1 vccd1 _11245_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_141_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09175__A _19693_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18841_ _19557_/CLK _18841_/D vssd1 vssd1 vccd1 vccd1 _18841_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09752__A2 _09741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ _11185_/A _11176_/B vssd1 vssd1 vccd1 vccd1 _11176_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10127_ _10127_/A _10127_/B vssd1 vssd1 vccd1 vccd1 _10127_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10993__S1 _10910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18772_ _19584_/CLK _18772_/D vssd1 vssd1 vccd1 vccd1 _18772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15984_ _15984_/A vssd1 vssd1 vccd1 vccd1 _18991_/D sky130_fd_sc_hd__clkbuf_1
X_17723_ _17723_/A vssd1 vssd1 vccd1 vccd1 _17772_/S sky130_fd_sc_hd__clkbuf_2
X_10058_ _18773_/Q _19002_/Q _18933_/Q _19231_/Q _09865_/A _10029_/A vssd1 vssd1 vccd1
+ vccd1 _10059_/B sky130_fd_sc_hd__mux4_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14935_ _18445_/Q _12632_/B _14981_/S vssd1 vssd1 vccd1 vccd1 _14935_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17654_ _17654_/A vssd1 vssd1 vccd1 vccd1 _19668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14866_ _16683_/A vssd1 vssd1 vccd1 vccd1 _16787_/A sky130_fd_sc_hd__buf_2
XFILLER_91_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16605_ _19258_/Q vssd1 vssd1 vccd1 vccd1 _16606_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__12686__D _13108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13817_ _13753_/X _13814_/Y _13816_/X vssd1 vssd1 vccd1 vccd1 _13817_/X sky130_fd_sc_hd__o21a_1
X_17585_ _17585_/A vssd1 vssd1 vccd1 vccd1 _19650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14797_ _15060_/B vssd1 vssd1 vccd1 vccd1 _15051_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_17_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19324_ _19581_/CLK _19324_/D vssd1 vssd1 vccd1 vccd1 _19324_/Q sky130_fd_sc_hd__dfxtp_1
X_16536_ _19225_/Q _15535_/X _16536_/S vssd1 vssd1 vccd1 vccd1 _16537_/A sky130_fd_sc_hd__mux2_1
X_13748_ _13746_/X _13747_/X _13877_/S vssd1 vssd1 vccd1 vccd1 _13748_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11170__S1 _09704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19255_ _19710_/CLK _19255_/D vssd1 vssd1 vccd1 vccd1 _19255_/Q sky130_fd_sc_hd__dfxtp_1
X_16467_ _16083_/X _19194_/Q _16475_/S vssd1 vssd1 vccd1 vccd1 _16468_/A sky130_fd_sc_hd__mux2_1
X_13679_ _12180_/A _14074_/B _13689_/S vssd1 vssd1 vccd1 vccd1 _13679_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18206_ _19856_/Q _18206_/B vssd1 vssd1 vccd1 vccd1 _18207_/B sky130_fd_sc_hd__xor2_1
X_15418_ _18753_/Q _15133_/X _15426_/S vssd1 vssd1 vccd1 vccd1 _15419_/A sky130_fd_sc_hd__mux2_1
X_19186_ _19634_/CLK _19186_/D vssd1 vssd1 vccd1 vccd1 _19186_/Q sky130_fd_sc_hd__dfxtp_1
X_16398_ _19164_/Q _15545_/X _16402_/S vssd1 vssd1 vccd1 vccd1 _16399_/A sky130_fd_sc_hd__mux2_1
X_18137_ _18140_/B _18140_/C _18126_/X vssd1 vssd1 vccd1 vccd1 _18137_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15349_ _18724_/Q _15149_/X _15351_/S vssd1 vssd1 vccd1 vccd1 _15350_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10050__A2 _10040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18068_ _18067_/B _18067_/C _19809_/Q vssd1 vssd1 vccd1 vccd1 _18069_/C sky130_fd_sc_hd__a21oi_1
XFILLER_117_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09910_ _09217_/X _09903_/X _09905_/X _09909_/X _09249_/X vssd1 vssd1 vccd1 vccd1
+ _09910_/X sky130_fd_sc_hd__a311o_4
X_17019_ _19414_/Q _16677_/X _17025_/S vssd1 vssd1 vccd1 vccd1 _17020_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12504__A _12504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09841_ _09841_/A vssd1 vssd1 vccd1 vccd1 _09843_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10433__S0 _09632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _09772_/A vssd1 vssd1 vccd1 vccd1 _09995_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15029__A0 _18453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13335__A _18371_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17241__S _17241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11066__A1 _10807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11161__S1 _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09206_ _19694_/Q vssd1 vssd1 vccd1 vccd1 _10827_/A sky130_fd_sc_hd__clkinv_2
XFILLER_33_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10026__C1 _09988_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09137_ _10960_/A vssd1 vssd1 vccd1 vccd1 _10969_/A sky130_fd_sc_hd__buf_2
XFILLER_120_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09431__A1 _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15504__A1 _15503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10672__S0 _10614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_135_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09719__C1 _09248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12414__A _18379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11030_ _10548_/A _11027_/X _11029_/X vssd1 vssd1 vccd1 vccd1 _11030_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17416__S _17424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _12982_/B _12982_/C _18308_/Q vssd1 vssd1 vccd1 vccd1 _12983_/B sky130_fd_sc_hd__a21oi_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10727__S1 _10726_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _16744_/A _17391_/A vssd1 vssd1 vccd1 vccd1 _15010_/A sky130_fd_sc_hd__or2_2
XFILLER_73_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ _11984_/A _11984_/D vssd1 vssd1 vccd1 vccd1 _11932_/X sky130_fd_sc_hd__or2_1
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14651_ _14654_/A _17775_/B vssd1 vssd1 vccd1 vccd1 _14652_/A sky130_fd_sc_hd__and2_1
XFILLER_33_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11863_ _11913_/A vssd1 vssd1 vccd1 vccd1 _14026_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13602_ _13597_/X _13600_/X _13757_/S vssd1 vssd1 vccd1 vccd1 _13602_/X sky130_fd_sc_hd__mux2_1
X_10814_ _18853_/Q _19311_/Q _11028_/S vssd1 vssd1 vccd1 vccd1 _10814_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11057__A1 _10797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17370_ _16816_/X _19555_/Q _17374_/S vssd1 vssd1 vccd1 vccd1 _17371_/A sky130_fd_sc_hd__mux2_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ _11794_/A _12095_/B vssd1 vssd1 vccd1 vccd1 _11794_/Y sky130_fd_sc_hd__nor2_1
X_14582_ _14582_/A _14582_/B vssd1 vssd1 vccd1 vccd1 _14582_/Y sky130_fd_sc_hd__nand2_1
X_16321_ _16083_/X _19130_/Q _16329_/S vssd1 vssd1 vccd1 vccd1 _16322_/A sky130_fd_sc_hd__mux2_1
X_10745_ _10752_/A _10745_/B vssd1 vssd1 vccd1 vccd1 _10745_/X sky130_fd_sc_hd__or2_1
X_13533_ _11551_/Y _14565_/A _13537_/A _13171_/A vssd1 vssd1 vccd1 vccd1 _13534_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_158_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16990__S _16990_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12006__A0 _12481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19040_ _19622_/CLK _19040_/D vssd1 vssd1 vccd1 vccd1 _19040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13464_ _18392_/Q _13245_/X _13464_/S vssd1 vssd1 vccd1 vccd1 _13465_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16252_ _16252_/A vssd1 vssd1 vccd1 vccd1 _19099_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16940__A0 _16771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10676_ _19691_/Q vssd1 vssd1 vccd1 vccd1 _10983_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_167_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10017__C1 _09988_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12415_ _18379_/Q _12414_/B _17693_/A vssd1 vssd1 vccd1 vccd1 _12415_/Y sky130_fd_sc_hd__o21ai_1
X_15203_ _16705_/A vssd1 vssd1 vccd1 vccd1 _15203_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13395_ _18263_/Q _12582_/A _12584_/A _19852_/Q vssd1 vssd1 vccd1 vccd1 _13395_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16183_ _16096_/X _19065_/Q _16183_/S vssd1 vssd1 vccd1 vccd1 _16184_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15134_ _15134_/A vssd1 vssd1 vccd1 vccd1 _15412_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12346_ _14580_/A _13525_/A _12345_/X _12501_/A vssd1 vssd1 vccd1 vccd1 _12347_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09973__A2 _09963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15065_ _16737_/A vssd1 vssd1 vccd1 vccd1 _16841_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14015__S _14032_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12277_ _14572_/A _12277_/B vssd1 vssd1 vccd1 vccd1 _12277_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14016_ _14016_/A vssd1 vssd1 vccd1 vccd1 _18433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output73_A _12511_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ _11229_/A _11227_/C _11227_/A vssd1 vssd1 vccd1 vccd1 _11228_/X sky130_fd_sc_hd__a21o_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15259__B1 _11822_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__S1 _10365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18824_ _19540_/CLK _18824_/D vssd1 vssd1 vccd1 vccd1 _18824_/Q sky130_fd_sc_hd__dfxtp_1
X_11159_ _10103_/A _11156_/X _11158_/X vssd1 vssd1 vccd1 vccd1 _11159_/X sky130_fd_sc_hd__a21o_1
XFILLER_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18755_ _19698_/CLK _18755_/D vssd1 vssd1 vccd1 vccd1 _18755_/Q sky130_fd_sc_hd__dfxtp_1
X_15967_ _15967_/A vssd1 vssd1 vccd1 vccd1 _18983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17706_ _17706_/A vssd1 vssd1 vccd1 vccd1 _19677_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16759__A0 _16758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14918_ _16800_/A vssd1 vssd1 vccd1 vccd1 _14918_/X sky130_fd_sc_hd__clkbuf_2
X_18686_ _19780_/CLK _18686_/D vssd1 vssd1 vccd1 vccd1 _18686_/Q sky130_fd_sc_hd__dfxtp_1
X_15898_ _14792_/X _18952_/Q _15902_/S vssd1 vssd1 vccd1 vccd1 _15899_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17637_ _19665_/Q _17636_/X _17653_/S vssd1 vssd1 vccd1 vccd1 _17638_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14849_ _14849_/A vssd1 vssd1 vccd1 vccd1 _18597_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12994__A _13034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16466__A _16488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17568_ _19643_/Q _16790_/A _17568_/S vssd1 vssd1 vccd1 vccd1 _17569_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19307_ _19691_/CLK _19307_/D vssd1 vssd1 vccd1 vccd1 _19307_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17184__A0 _18439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16519_ _19217_/Q _15510_/X _16525_/S vssd1 vssd1 vccd1 vccd1 _16520_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17499_ _19612_/Q _16689_/X _17507_/S vssd1 vssd1 vccd1 vccd1 _17500_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19238_ _19643_/CLK _19238_/D vssd1 vssd1 vccd1 vccd1 _19238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16931__A0 _16758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10507__B_N _12478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09949__C1 _09395_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19169_ _19718_/CLK _19169_/D vssd1 vssd1 vccd1 vccd1 _19169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16405__S _16413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10654__S0 _10836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10406__S0 _09673_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10957__S1 _10910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12720__B2 _19481_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09824_ _09952_/S vssd1 vssd1 vccd1 vccd1 _09874_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_150_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09755_ _09755_/A _09901_/A vssd1 vssd1 vccd1 vccd1 _11224_/A sky130_fd_sc_hd__nor2_1
XFILLER_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09686_ _18453_/Q _09309_/A _09429_/A _09685_/X vssd1 vssd1 vccd1 vccd1 _12501_/A
+ sky130_fd_sc_hd__o2bb2a_4
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15280__A _15337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_61_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12409__A _19757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10798__B1 _10944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17714__A2 _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10530_ _10566_/A _10530_/B vssd1 vssd1 vccd1 vccd1 _10530_/X sky130_fd_sc_hd__or2_1
XFILLER_167_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10461_ _10461_/A _12480_/A vssd1 vssd1 vccd1 vccd1 _10462_/B sky130_fd_sc_hd__or2_1
XFILLER_108_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12200_ _12196_/X _12198_/X _12199_/Y _11801_/X vssd1 vssd1 vccd1 vccd1 _12200_/X
+ sky130_fd_sc_hd__a31o_1
X_13180_ _19828_/Q _12736_/A _13175_/X _13177_/X _13179_/X vssd1 vssd1 vccd1 vccd1
+ _13181_/B sky130_fd_sc_hd__a2111o_4
X_10392_ _10392_/A vssd1 vssd1 vccd1 vccd1 _10442_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12131_ _12131_/A _12131_/B _12131_/C _12131_/D vssd1 vssd1 vccd1 vccd1 _12132_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__12144__A _19745_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14161__A0 _18442_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12062_ _12063_/A _13603_/A vssd1 vssd1 vccd1 vccd1 _12064_/A sky130_fd_sc_hd__and2_1
XFILLER_151_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11013_ _19502_/Q _19116_/Q _19566_/Q _18722_/Q _09336_/A _10940_/X vssd1 vssd1 vccd1
+ vccd1 _11014_/B sky130_fd_sc_hd__mux4_2
XFILLER_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16870_ _16870_/A vssd1 vssd1 vccd1 vccd1 _19348_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15821_ _15878_/S vssd1 vssd1 vccd1 vccd1 _15830_/S sky130_fd_sc_hd__buf_2
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18540_ _18548_/CLK _18540_/D vssd1 vssd1 vccd1 vccd1 _18540_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _14782_/X _18887_/Q _15758_/S vssd1 vssd1 vccd1 vccd1 _15753_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _18303_/Q vssd1 vssd1 vccd1 vccd1 _12972_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14703_ _14703_/A vssd1 vssd1 vccd1 vccd1 _14703_/X sky130_fd_sc_hd__buf_2
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ _14059_/B _11915_/B vssd1 vssd1 vccd1 vccd1 _11918_/A sky130_fd_sc_hd__xnor2_1
X_18471_ _18471_/CLK _18471_/D vssd1 vssd1 vccd1 vccd1 _18471_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15683_ _15683_/A vssd1 vssd1 vccd1 vccd1 _18856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12895_ _18278_/Q _18277_/Q _12895_/C _12895_/D vssd1 vssd1 vccd1 vccd1 _12933_/C
+ sky130_fd_sc_hd__and4_2
XFILLER_166_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17422_ _16787_/X _19578_/Q _17424_/S vssd1 vssd1 vccd1 vccd1 _17423_/A sky130_fd_sc_hd__mux2_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ _18565_/Q _14633_/X _14622_/X input36/X vssd1 vssd1 vccd1 vccd1 _14635_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _11846_/A _11846_/B vssd1 vssd1 vccd1 vccd1 _11846_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13422__B _13422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17353_ _17353_/A vssd1 vssd1 vccd1 vccd1 _19547_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ _14565_/A vssd1 vssd1 vccd1 vccd1 _14580_/B sky130_fd_sc_hd__clkbuf_1
X_11777_ _11733_/B _14036_/S _11970_/A vssd1 vssd1 vccd1 vccd1 _11778_/B sky130_fd_sc_hd__a21o_1
XFILLER_60_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _16304_/A vssd1 vssd1 vccd1 vccd1 _19122_/D sky130_fd_sc_hd__clkbuf_1
X_13516_ _14601_/A _13516_/B vssd1 vssd1 vccd1 vccd1 _13563_/A sky130_fd_sc_hd__and2_1
X_10728_ _10728_/A vssd1 vssd1 vccd1 vccd1 _10728_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_158_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17284_ _17284_/A vssd1 vssd1 vccd1 vccd1 _19516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14496_ _18518_/Q _19756_/Q _14498_/S vssd1 vssd1 vccd1 vccd1 _14497_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13727__B1 _13723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19023_ _19713_/CLK _19023_/D vssd1 vssd1 vccd1 vccd1 _19023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16235_ _16064_/X _19092_/Q _16235_/S vssd1 vssd1 vccd1 vccd1 _16236_/A sky130_fd_sc_hd__mux2_1
X_13447_ _18384_/Q _13149_/X _13453_/S vssd1 vssd1 vccd1 vccd1 _13448_/A sky130_fd_sc_hd__mux2_1
X_10659_ _18434_/Q _09307_/A _09428_/A _10658_/X vssd1 vssd1 vccd1 vccd1 _12473_/A
+ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__14534__A _17892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09628__A _11200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13378_ _13354_/X _13376_/X _13377_/X _13350_/X vssd1 vssd1 vccd1 vccd1 _18376_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16166_ _16071_/X _19057_/Q _16172_/S vssd1 vssd1 vccd1 vccd1 _16167_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12950__A1 _18293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15117_ _18638_/Q _15116_/X _15111_/X _11139_/A vssd1 vssd1 vccd1 vccd1 _18638_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12329_ _11222_/A _18516_/Q _12423_/S vssd1 vssd1 vccd1 vccd1 _12355_/A sky130_fd_sc_hd__mux2_8
XFILLER_173_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16097_ _16096_/X _19033_/Q _16097_/S vssd1 vssd1 vccd1 vccd1 _16098_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15048_ _17765_/A _15049_/B vssd1 vssd1 vccd1 vccd1 _15048_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17056__S _17058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11893__A _11940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19856_ _19856_/CLK _19856_/D vssd1 vssd1 vccd1 vccd1 _19856_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_122_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09363__A _09826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18807_ _19587_/CLK _18807_/D vssd1 vssd1 vccd1 vccd1 _18807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19787_ _19795_/CLK _19787_/D vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dfxtp_1
XFILLER_84_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16999_ _19405_/Q _16648_/X _17003_/S vssd1 vssd1 vccd1 vccd1 _17000_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09540_ _09554_/A vssd1 vssd1 vccd1 vccd1 _10306_/A sky130_fd_sc_hd__buf_4
XFILLER_77_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18738_ _19613_/CLK _18738_/D vssd1 vssd1 vccd1 vccd1 _18738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10302__A _10313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09471_ _09275_/A _09461_/X _09470_/X _09282_/A _18456_/Q vssd1 vssd1 vccd1 vccd1
+ _11202_/A sky130_fd_sc_hd__a32o_4
X_18669_ _19714_/CLK _18669_/D vssd1 vssd1 vccd1 vccd1 _18669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17157__A0 _18431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16135__S _16135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09538__A _09538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10183__S _11188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12899__A _18279_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09807_ _10055_/S vssd1 vssd1 vccd1 vccd1 _09808_/A sky130_fd_sc_hd__buf_2
XFILLER_115_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14446__A1 _19733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10180__A1 _09414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09738_ _19429_/Q _19205_/Q _19722_/Q _19173_/Q _09729_/S _09728_/A vssd1 vssd1 vccd1
+ vccd1 _09738_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10212__A _10212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17396__A0 _16749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _09412_/A _09659_/Y _09661_/Y _09666_/Y _09668_/Y vssd1 vssd1 vccd1 vccd1
+ _09669_/X sky130_fd_sc_hd__o32a_1
XANTENNA__15214__S _15217_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11700_ _11746_/A _11700_/B vssd1 vssd1 vccd1 vccd1 _11703_/B sky130_fd_sc_hd__or2_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13523__A _14584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12680_ _19859_/Q _12582_/X _12584_/X _19827_/Q vssd1 vssd1 vccd1 vccd1 _12680_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10483__A2 _10473_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14749__A2 _12683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11997_/A _11630_/X _17855_/C _19729_/Q vssd1 vssd1 vccd1 vccd1 _17857_/B
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13421__A2 _12665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11562_ _12017_/B vssd1 vssd1 vccd1 vccd1 _12412_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14350_ _14350_/A vssd1 vssd1 vccd1 vccd1 _18461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13301_ _19484_/Q _13203_/A _13205_/A _18398_/Q vssd1 vssd1 vccd1 vccd1 _13301_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10513_ _10227_/A _10508_/X _10510_/X _10512_/X vssd1 vssd1 vccd1 vccd1 _10513_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14281_ _12333_/X _14102_/X _14280_/X vssd1 vssd1 vccd1 vccd1 _14281_/X sky130_fd_sc_hd__a21bo_1
X_11493_ _11513_/A _11514_/A _13524_/C vssd1 vssd1 vccd1 vccd1 _11519_/C sky130_fd_sc_hd__or3_1
XFILLER_155_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16020_ _16020_/A vssd1 vssd1 vccd1 vccd1 _19007_/D sky130_fd_sc_hd__clkbuf_1
X_13232_ _17781_/A vssd1 vssd1 vccd1 vccd1 _13232_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_input72_A reset vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10444_ _10438_/A _10443_/X _09411_/A vssd1 vssd1 vccd1 vccd1 _10444_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09484__S0 _10389_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13163_ _18621_/Q _13163_/B vssd1 vssd1 vccd1 vccd1 _13163_/X sky130_fd_sc_hd__or2_1
XFILLER_152_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10375_ _10428_/A _10375_/B vssd1 vssd1 vccd1 vccd1 _10375_/X sky130_fd_sc_hd__or2_1
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12114_ _12114_/A _12114_/B vssd1 vssd1 vccd1 vccd1 _14163_/A sky130_fd_sc_hd__xnor2_4
XFILLER_97_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13094_ input67/X _13104_/B vssd1 vssd1 vccd1 vccd1 _13094_/X sky130_fd_sc_hd__or2_1
X_17971_ _19775_/Q _19774_/Q _17971_/C vssd1 vssd1 vccd1 vccd1 _17973_/B sky130_fd_sc_hd__and3_1
XFILLER_97_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19710_ _19710_/CLK _19710_/D vssd1 vssd1 vccd1 vccd1 _19710_/Q sky130_fd_sc_hd__dfxtp_1
X_12045_ _12041_/A _12044_/X _12119_/S vssd1 vssd1 vccd1 vccd1 _12045_/X sky130_fd_sc_hd__mux2_1
X_16922_ _16990_/S vssd1 vssd1 vccd1 vccd1 _16931_/S sky130_fd_sc_hd__buf_2
XANTENNA__09787__S1 _09763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12602__A _12602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19641_ _19710_/CLK _19641_/D vssd1 vssd1 vccd1 vccd1 _19641_/Q sky130_fd_sc_hd__dfxtp_1
X_16853_ _16853_/A vssd1 vssd1 vccd1 vccd1 _19340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14437__A1 _19729_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10171__B2 _18444_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15804_ _15066_/X _18911_/Q _15806_/S vssd1 vssd1 vccd1 vccd1 _15805_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19572_ _19702_/CLK _19572_/D vssd1 vssd1 vccd1 vccd1 _19572_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12448__B1 _13702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16784_ _16784_/A vssd1 vssd1 vccd1 vccd1 _16784_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_92_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13996_ _13996_/A _13996_/B vssd1 vssd1 vccd1 vccd1 _13996_/X sky130_fd_sc_hd__and2_1
XFILLER_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18523_ _18564_/CLK _18523_/D vssd1 vssd1 vccd1 vccd1 _18523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15735_ _15735_/A vssd1 vssd1 vccd1 vccd1 _18880_/D sky130_fd_sc_hd__clkbuf_1
X_12947_ _12983_/A _12947_/B _12952_/C vssd1 vssd1 vccd1 vccd1 _18292_/D sky130_fd_sc_hd__nor3_1
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09864__B2 _18451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ _18632_/CLK _18454_/D vssd1 vssd1 vccd1 vccd1 _18454_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15666_ _15734_/S vssd1 vssd1 vccd1 vccd1 _15675_/S sky130_fd_sc_hd__buf_2
X_12878_ _18272_/Q _12874_/C _12877_/Y vssd1 vssd1 vccd1 vccd1 _18272_/D sky130_fd_sc_hd__o21a_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _16761_/X _19570_/Q _17413_/S vssd1 vssd1 vccd1 vccd1 _17406_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13152__B _18621_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14617_ input62/X _14593_/X _14597_/X _14524_/A vssd1 vssd1 vccd1 vccd1 _14618_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18385_ _19780_/CLK _18385_/D vssd1 vssd1 vccd1 vccd1 _18385_/Q sky130_fd_sc_hd__dfxtp_1
X_11829_ _15262_/A _11828_/X _11801_/A vssd1 vssd1 vccd1 vccd1 _11829_/X sky130_fd_sc_hd__a21o_1
XFILLER_159_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15597_ _18818_/Q _15494_/X _15603_/S vssd1 vssd1 vccd1 vccd1 _15598_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16744__A _16744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17336_ _17336_/A vssd1 vssd1 vccd1 vccd1 _19539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09711__S1 _10080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14548_ _14585_/A vssd1 vssd1 vccd1 vccd1 _14548_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17267_ _19509_/Q _16667_/X _17269_/S vssd1 vssd1 vccd1 vccd1 _17268_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14479_ _18510_/Q _19748_/Q _14487_/S vssd1 vssd1 vccd1 vccd1 _14480_/A sky130_fd_sc_hd__mux2_1
X_19006_ _19589_/CLK _19006_/D vssd1 vssd1 vccd1 vccd1 _19006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09358__A _10329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16218_ _16039_/X _19084_/Q _16224_/S vssd1 vssd1 vccd1 vccd1 _16219_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17198_ _18443_/Q _12598_/B _17201_/S vssd1 vssd1 vccd1 vccd1 _17198_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15794__S _15802_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16149_ _16149_/A vssd1 vssd1 vccd1 vccd1 _19049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14676__A1 _14575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14676__B2 input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15095__A _15095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13608__A _13608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12512__A _18417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19839_ _19851_/CLK _19839_/D vssd1 vssd1 vccd1 vccd1 _19839_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15625__A0 _18831_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17514__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09523_ _18847_/Q _19401_/Q _19563_/Q _18815_/Q _11110_/S _09587_/A vssd1 vssd1 vccd1
+ vccd1 _09524_/B sky130_fd_sc_hd__mux4_1
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15034__S _15056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09454_ _09454_/A vssd1 vssd1 vccd1 vccd1 _09463_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09385_ _09385_/A vssd1 vssd1 vccd1 vccd1 _09814_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09607__A1 _09414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09466__S0 _10465_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10160_ _09996_/A _10157_/X _10159_/X _09230_/A vssd1 vssd1 vccd1 vccd1 _10160_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11025__S0 _10919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ _10107_/A _10090_/X _10007_/A vssd1 vssd1 vccd1 vccd1 _10091_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11433__A1_N _12555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12422__A _14324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14419__A1 _18517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17424__S _17424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13850_ _13846_/Y _13946_/A _13995_/S vssd1 vssd1 vccd1 vccd1 _13850_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15092__A1 _10834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12801_ _13042_/A vssd1 vssd1 vccd1 vccd1 _18173_/A sky130_fd_sc_hd__buf_2
XFILLER_142_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13781_ _14019_/S vssd1 vssd1 vccd1 vccd1 _14122_/S sky130_fd_sc_hd__clkbuf_2
X_10993_ _19630_/Q _19047_/Q _19084_/Q _18690_/Q _10909_/X _10910_/X vssd1 vssd1 vccd1
+ vccd1 _10993_/X sky130_fd_sc_hd__mux4_2
XANTENNA__12795__C _18214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15520_ _18794_/Q _15519_/X _15520_/S vssd1 vssd1 vccd1 vccd1 _15521_/A sky130_fd_sc_hd__mux2_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12732_ _18299_/Q _12810_/A vssd1 vssd1 vccd1 vccd1 _12732_/X sky130_fd_sc_hd__or2_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09941__S1 _09881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _18768_/Q _15187_/X _15459_/S vssd1 vssd1 vccd1 vccd1 _15452_/A sky130_fd_sc_hd__mux2_1
X_12663_ _13178_/A vssd1 vssd1 vccd1 vccd1 _12663_/X sky130_fd_sc_hd__buf_2
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14783__S _14822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14402_ _14402_/A vssd1 vssd1 vccd1 vccd1 _18479_/D sky130_fd_sc_hd__clkbuf_1
X_18170_ _18170_/A vssd1 vssd1 vccd1 vccd1 _18170_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11614_ _18562_/Q _11371_/Y _11835_/S _12277_/B _11613_/X vssd1 vssd1 vccd1 vccd1
+ _11614_/X sky130_fd_sc_hd__o2111a_2
XFILLER_168_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15382_ _18739_/Q _15197_/X _15384_/S vssd1 vssd1 vccd1 vccd1 _15383_/A sky130_fd_sc_hd__mux2_1
X_12594_ _18636_/Q _12594_/B vssd1 vssd1 vccd1 vccd1 _12594_/X sky130_fd_sc_hd__or2_1
X_17121_ _17121_/A vssd1 vssd1 vccd1 vccd1 _17130_/S sky130_fd_sc_hd__buf_4
X_14333_ _13937_/X _12446_/B _14088_/A _14332_/X vssd1 vssd1 vccd1 vccd1 _14333_/X
+ sky130_fd_sc_hd__o211a_1
X_11545_ _11545_/A vssd1 vssd1 vccd1 vccd1 _19080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13158__B2 _19661_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17052_ _19429_/Q _16725_/X _17058_/S vssd1 vssd1 vccd1 vccd1 _17053_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09178__A _10996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14264_ _13975_/X _14261_/Y _14263_/X _13721_/X vssd1 vssd1 vccd1 vccd1 _14264_/X
+ sky130_fd_sc_hd__a211o_1
X_11476_ _13583_/B _11476_/B vssd1 vssd1 vccd1 vccd1 _13570_/D sky130_fd_sc_hd__nor2_2
XFILLER_143_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16003_ _14929_/X _19000_/Q _16005_/S vssd1 vssd1 vccd1 vccd1 _16004_/A sky130_fd_sc_hd__mux2_1
X_13215_ _13215_/A _13246_/B vssd1 vssd1 vccd1 vccd1 _13215_/X sky130_fd_sc_hd__or2_1
X_10427_ _19513_/Q _19127_/Q _19577_/Q _18733_/Q _11087_/S _10368_/X vssd1 vssd1 vccd1
+ vccd1 _10428_/B sky130_fd_sc_hd__mux4_1
XFILLER_136_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14195_ _13971_/X _14086_/X _14194_/X vssd1 vssd1 vccd1 vccd1 _14195_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_183_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13146_ _12972_/B _13130_/X _12664_/A _18023_/B _13145_/X vssd1 vssd1 vccd1 vccd1
+ _13146_/X sky130_fd_sc_hd__a221o_1
X_10358_ _10866_/A vssd1 vssd1 vccd1 vccd1 _10752_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17954_ _19769_/Q _17954_/B _17954_/C vssd1 vssd1 vccd1 vccd1 _17955_/C sky130_fd_sc_hd__and3_1
XFILLER_151_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13077_ _19799_/Q vssd1 vssd1 vccd1 vccd1 _18043_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _19645_/Q _19062_/Q _19099_/Q _18705_/Q _09675_/S _10239_/X vssd1 vssd1 vccd1
+ vccd1 _10289_/X sky130_fd_sc_hd__mux4_2
XFILLER_140_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16905_ _19364_/Q _16721_/X _16913_/S vssd1 vssd1 vccd1 vccd1 _16906_/A sky130_fd_sc_hd__mux2_1
X_12028_ _12155_/A _12028_/B vssd1 vssd1 vccd1 vccd1 _12131_/A sky130_fd_sc_hd__nand2_1
XFILLER_78_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17885_ _17885_/A vssd1 vssd1 vccd1 vccd1 _19743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16836_ _16835_/X _19335_/Q _16839_/S vssd1 vssd1 vccd1 vccd1 _16837_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19624_ _19624_/CLK _19624_/D vssd1 vssd1 vccd1 vccd1 _19624_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11892__A1 _12474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19710_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11892__B2 _11513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19555_ _19555_/CLK _19555_/D vssd1 vssd1 vccd1 vccd1 _19555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16767_ _16767_/A vssd1 vssd1 vccd1 vccd1 _19313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09837__A1 _09320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13979_ _14040_/A vssd1 vssd1 vccd1 vccd1 _13979_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14830__A1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13163__A _18621_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18506_ _18506_/CLK _18506_/D vssd1 vssd1 vccd1 vccd1 _18506_/Q sky130_fd_sc_hd__dfxtp_1
X_15718_ _15718_/A vssd1 vssd1 vccd1 vccd1 _18872_/D sky130_fd_sc_hd__clkbuf_1
X_19486_ _19488_/CLK _19486_/D vssd1 vssd1 vccd1 vccd1 _19486_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09932__S1 _09869_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16698_ _16698_/A vssd1 vssd1 vccd1 vccd1 _19292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15789__S _15791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18437_ _18818_/CLK _18437_/D vssd1 vssd1 vccd1 vccd1 _18437_/Q sky130_fd_sc_hd__dfxtp_4
X_15649_ _15649_/A vssd1 vssd1 vccd1 vccd1 _15658_/S sky130_fd_sc_hd__buf_4
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09170_ _09170_/A vssd1 vssd1 vccd1 vccd1 _09171_/A sky130_fd_sc_hd__clkbuf_4
X_18368_ _18402_/CLK _18368_/D vssd1 vssd1 vccd1 vccd1 _18368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17319_ _17783_/A _17319_/B vssd1 vssd1 vccd1 vccd1 _17376_/A sky130_fd_sc_hd__nand2_4
XFILLER_147_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18299_ _19856_/CLK _18299_/D vssd1 vssd1 vccd1 vccd1 _18299_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09470__C1 _09246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13149__B2 _18620_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14897__A1 _12554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11130__B _12481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10058__S1 _10029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16413__S _16413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09999__S1 _09763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14722__A _15077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10383__B2 _18440_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09620__S0 _09344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13085__B1 _12602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09506_ _10400_/A _09506_/B vssd1 vssd1 vccd1 vccd1 _09506_/Y sky130_fd_sc_hd__nor2_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09437_ _10982_/S vssd1 vssd1 vccd1 vccd1 _10733_/S sky130_fd_sc_hd__buf_2
XFILLER_53_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09368_ _09368_/A vssd1 vssd1 vccd1 vccd1 _09368_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09299_ _18532_/Q vssd1 vssd1 vccd1 vccd1 _15412_/B sky130_fd_sc_hd__inv_2
XANTENNA__09461__C1 _10373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _18584_/Q _18583_/Q _18582_/Q _18581_/Q vssd1 vssd1 vccd1 vccd1 _11344_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17927__B _19760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12136__B _13596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11261_ _11261_/A _11261_/B _11261_/C _11260_/X vssd1 vssd1 vccd1 vccd1 _11261_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_137_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16323__S _16329_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13000_ _13003_/B _13003_/C _12922_/X vssd1 vssd1 vccd1 vccd1 _13000_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_107_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10212_ _10212_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10212_/X sky130_fd_sc_hd__or2_1
X_11192_ _19431_/Q _19207_/Q _19724_/Q _19175_/Q _11186_/S _10329_/A vssd1 vssd1 vccd1
+ vccd1 _11192_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11975__B _12011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10143_ _18836_/Q _19390_/Q _19552_/Q _18804_/Q _10125_/X _09867_/A vssd1 vssd1 vccd1
+ vccd1 _10144_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12152__A _19746_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input35_A io_ibus_inst[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ _10074_/A _10074_/B vssd1 vssd1 vccd1 vccd1 _10074_/X sky130_fd_sc_hd__or2_1
X_14951_ _16809_/A vssd1 vssd1 vccd1 vccd1 _14951_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09611__S0 _10131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13902_ _14285_/A _14103_/A vssd1 vssd1 vccd1 vccd1 _13902_/X sky130_fd_sc_hd__or2_1
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17670_ _12727_/X _17669_/Y _17686_/S vssd1 vssd1 vccd1 vccd1 _17670_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10221__S1 _09602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14882_ input7/X _14801_/A _14804_/A vssd1 vssd1 vccd1 vccd1 _14887_/A sky130_fd_sc_hd__a21o_1
XFILLER_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16621_ _19266_/Q vssd1 vssd1 vccd1 vccd1 _16622_/A sky130_fd_sc_hd__clkbuf_1
X_13833_ _13880_/S _13833_/B vssd1 vssd1 vccd1 vccd1 _13833_/X sky130_fd_sc_hd__or2_1
XFILLER_29_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19340_ _19598_/CLK _19340_/D vssd1 vssd1 vccd1 vccd1 _19340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16552_ _19232_/Q _15558_/X _16558_/S vssd1 vssd1 vccd1 vccd1 _16553_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13764_ _13600_/X _13621_/X _13768_/S vssd1 vssd1 vccd1 vccd1 _13764_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10400__A _10400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _09208_/A _10973_/Y _10975_/Y _09243_/A vssd1 vssd1 vccd1 vccd1 _10976_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_15_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15503_ _16758_/A vssd1 vssd1 vccd1 vccd1 _15503_/X sky130_fd_sc_hd__clkbuf_2
X_12715_ _12715_/A _12715_/B vssd1 vssd1 vccd1 vccd1 _13516_/B sky130_fd_sc_hd__nand2_1
X_19271_ _19271_/CLK _19271_/D vssd1 vssd1 vccd1 vccd1 _19271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16483_ _16483_/A vssd1 vssd1 vccd1 vccd1 _19201_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17762__A0 _13412_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13695_ _14019_/S vssd1 vssd1 vccd1 vccd1 _14086_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__14807__A _16667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18222_ _19862_/Q _19861_/Q _18222_/C vssd1 vssd1 vccd1 vccd1 _18223_/B sky130_fd_sc_hd__and3_1
XANTENNA__15402__S _15406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15434_ _15434_/A vssd1 vssd1 vccd1 vccd1 _18760_/D sky130_fd_sc_hd__clkbuf_1
X_12646_ _18343_/Q _15242_/A _13418_/S _19489_/Q _12645_/X vssd1 vssd1 vccd1 vccd1
+ _12646_/X sky130_fd_sc_hd__a221o_1
XFILLER_129_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18153_ _19838_/Q _18156_/C _18126_/X vssd1 vssd1 vccd1 vccd1 _18153_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15365_ _18731_/Q _15171_/X _15373_/S vssd1 vssd1 vccd1 vccd1 _15366_/A sky130_fd_sc_hd__mux2_1
X_12577_ _13297_/A vssd1 vssd1 vccd1 vccd1 _12577_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_157_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17104_ _16800_/X _19452_/Q _17108_/S vssd1 vssd1 vccd1 vccd1 _17105_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ _13823_/X _13855_/Y _14315_/X _13871_/X vssd1 vssd1 vccd1 vccd1 _14316_/X
+ sky130_fd_sc_hd__a211o_1
X_18084_ _18086_/B _18086_/C _18083_/Y vssd1 vssd1 vccd1 vccd1 _19814_/D sky130_fd_sc_hd__o21a_1
X_11528_ _11528_/A _11528_/B vssd1 vssd1 vccd1 vccd1 _11599_/B sky130_fd_sc_hd__or2_1
X_15296_ _18701_/Q _15178_/X _15300_/S vssd1 vssd1 vccd1 vccd1 _15297_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12339__C1 _12193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17035_ _17035_/A vssd1 vssd1 vccd1 vccd1 _19421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13000__B1 _12922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14247_ _18449_/Q _14246_/X _14306_/S vssd1 vssd1 vccd1 vccd1 _14248_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11459_ _15093_/S vssd1 vssd1 vccd1 vccd1 _11460_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09636__A _10349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ _14178_/A _14178_/B vssd1 vssd1 vccd1 vccd1 _14178_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_140_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _18506_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__15828__A0 _14808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14261__B _14265_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09850__S0 _09914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13129_ _18684_/Q _12671_/X _13125_/X _13128_/X vssd1 vssd1 vccd1 vccd1 _13129_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_124_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18986_ _19601_/CLK _18986_/D vssd1 vssd1 vccd1 vccd1 _18986_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13303__A1 _19674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17937_ _17946_/D vssd1 vssd1 vccd1 vccd1 _17944_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10117__A1 _09979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12997__A _12997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17868_ _17874_/A _17868_/B vssd1 vssd1 vccd1 vccd1 _17869_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_155_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19700_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19607_ _19706_/CLK _19607_/D vssd1 vssd1 vccd1 vccd1 _19607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16819_ _16819_/A vssd1 vssd1 vccd1 vccd1 _16819_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17799_ _15159_/X _19702_/Q _17805_/S vssd1 vssd1 vccd1 vccd1 _17800_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11406__A _13130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19538_ _19539_/CLK _19538_/D vssd1 vssd1 vccd1 vccd1 _19538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19469_ _19472_/CLK _19469_/D vssd1 vssd1 vccd1 vccd1 _19469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09222_ _19694_/Q vssd1 vssd1 vccd1 vccd1 _09223_/A sky130_fd_sc_hd__buf_2
XFILLER_10_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ _10605_/S vssd1 vssd1 vccd1 vccd1 _10604_/S sky130_fd_sc_hd__buf_2
XFILLER_30_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11141__A _12491_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09994__B1 _10007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09084_ _18559_/Q vssd1 vssd1 vccd1 vccd1 _11321_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_163_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_108_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19753_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15267__B _17535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09986_ _10022_/A _09986_/B vssd1 vssd1 vccd1 vccd1 _09986_/X sky130_fd_sc_hd__or2_1
XFILLER_88_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12700__A _12766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15047__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10830_ _10830_/A _10830_/B vssd1 vssd1 vccd1 vccd1 _10830_/X sky130_fd_sc_hd__or2_1
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_131_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10761_ _18823_/Q _19377_/Q _19539_/Q _18791_/Q _10836_/A _09482_/A vssd1 vssd1 vccd1
+ vccd1 _10762_/B sky130_fd_sc_hd__mux4_2
XANTENNA__16318__S _16318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12500_ _12500_/A _12503_/B vssd1 vssd1 vccd1 vccd1 _12500_/Y sky130_fd_sc_hd__nor2_1
X_13480_ _18399_/Q _12559_/X _13486_/S vssd1 vssd1 vccd1 vccd1 _13481_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10692_ _11056_/A vssd1 vssd1 vccd1 vccd1 _10701_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12431_ _12431_/A _12431_/B vssd1 vssd1 vccd1 vccd1 _14319_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__12033__A1 _18504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15150_ _18654_/Q _15149_/X _15153_/S vssd1 vssd1 vccd1 vccd1 _15151_/A sky130_fd_sc_hd__mux2_1
X_12362_ _12362_/A _12386_/B vssd1 vssd1 vccd1 vccd1 _12362_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14101_ _18438_/Q _11460_/X _14100_/X vssd1 vssd1 vccd1 vccd1 _18438_/D sky130_fd_sc_hd__o21a_1
XFILLER_165_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11313_ _11365_/B _11339_/B _12471_/B _11313_/D vssd1 vssd1 vccd1 vccd1 _11599_/A
+ sky130_fd_sc_hd__or4_2
X_12293_ _12293_/A _12335_/C vssd1 vssd1 vccd1 vccd1 _12293_/Y sky130_fd_sc_hd__nor2_1
X_15081_ _18619_/Q _15080_/X _15087_/S vssd1 vssd1 vccd1 vccd1 _15082_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16053__S _16065_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14730__A0 _14729_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09456__A _10622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14032_ _18434_/Q _14031_/Y _14032_/S vssd1 vssd1 vccd1 vccd1 _14033_/A sky130_fd_sc_hd__mux2_1
X_11244_ _11244_/A _11244_/B vssd1 vssd1 vccd1 vccd1 _11247_/B sky130_fd_sc_hd__nor2_1
XFILLER_153_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13533__B2 _13171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11544__A0 _11542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16988__S _16990_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18840_ _19556_/CLK _18840_/D vssd1 vssd1 vccd1 vccd1 _18840_/Q sky130_fd_sc_hd__dfxtp_1
X_11175_ _19625_/Q _19463_/Q _18909_/Q _18679_/Q _10129_/S _09736_/A vssd1 vssd1 vccd1
+ vccd1 _11176_/B sky130_fd_sc_hd__mux4_1
XFILLER_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09752__A3 _09750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_72_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19295_/CLK sky130_fd_sc_hd__clkbuf_16
X_10126_ _19262_/Q _19033_/Q _18964_/Q _19358_/Q _10125_/X _09595_/A vssd1 vssd1 vccd1
+ vccd1 _10127_/B sky130_fd_sc_hd__mux4_1
XFILLER_121_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18771_ _19714_/CLK _18771_/D vssd1 vssd1 vccd1 vccd1 _18771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15983_ _14821_/X _18991_/Q _15983_/S vssd1 vssd1 vccd1 vccd1 _15984_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17722_ _17728_/B _17721_/Y _17711_/X vssd1 vssd1 vccd1 vccd1 _17722_/Y sky130_fd_sc_hd__a21oi_1
X_10057_ _10064_/A _10052_/X _10054_/X _10056_/X vssd1 vssd1 vccd1 vccd1 _10057_/X
+ sky130_fd_sc_hd__o22a_1
X_14934_ _14969_/A _14955_/C _14934_/C vssd1 vssd1 vccd1 vccd1 _14934_/X sky130_fd_sc_hd__or3_2
XFILLER_75_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17653_ _19668_/Q _17652_/X _17653_/S vssd1 vssd1 vccd1 vccd1 _17654_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14865_ _14811_/X _14860_/X _14863_/X _14864_/X vssd1 vssd1 vccd1 vccd1 _16683_/A
+ sky130_fd_sc_hd__o31a_4
XFILLER_63_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_87_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19790_/CLK sky130_fd_sc_hd__clkbuf_16
X_16604_ _16604_/A vssd1 vssd1 vccd1 vccd1 _19257_/D sky130_fd_sc_hd__clkbuf_1
X_13816_ _13816_/A vssd1 vssd1 vccd1 vccd1 _13816_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17584_ _19650_/Q _16813_/A _17590_/S vssd1 vssd1 vccd1 vccd1 _17585_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14796_ _18466_/Q _14796_/B vssd1 vssd1 vccd1 vccd1 _14827_/C sky130_fd_sc_hd__and2_1
XFILLER_44_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19323_ _19581_/CLK _19323_/D vssd1 vssd1 vccd1 vccd1 _19323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16535_ _16535_/A vssd1 vssd1 vccd1 vccd1 _19224_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17735__A0 _19682_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13747_ _13672_/X _13666_/X _13747_/S vssd1 vssd1 vccd1 vccd1 _13747_/X sky130_fd_sc_hd__mux2_1
X_10959_ _10959_/A vssd1 vssd1 vccd1 vccd1 _10959_/X sky130_fd_sc_hd__buf_4
XANTENNA__14537__A _15412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19254_ _19414_/CLK _19254_/D vssd1 vssd1 vccd1 vccd1 _19254_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_10_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19723_/CLK sky130_fd_sc_hd__clkbuf_16
X_16466_ _16488_/A vssd1 vssd1 vccd1 vccd1 _16475_/S sky130_fd_sc_hd__buf_2
X_13678_ _13623_/Y _14057_/B _13685_/S vssd1 vssd1 vccd1 vccd1 _13678_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_opt_3_0_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18205_ _18205_/A _18205_/B vssd1 vssd1 vccd1 vccd1 _18206_/B sky130_fd_sc_hd__nand2_1
X_15417_ _15485_/S vssd1 vssd1 vccd1 vccd1 _15426_/S sky130_fd_sc_hd__clkbuf_4
X_12629_ _19779_/Q _12627_/X _12629_/S vssd1 vssd1 vccd1 vccd1 _12629_/X sky130_fd_sc_hd__mux2_1
X_19185_ _19635_/CLK _19185_/D vssd1 vssd1 vccd1 vccd1 _19185_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13221__B1 _12742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12057__A _12057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16397_ _16397_/A vssd1 vssd1 vccd1 vccd1 _19163_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18136_ _19831_/Q _18132_/C _18135_/Y vssd1 vssd1 vccd1 vccd1 _19831_/D sky130_fd_sc_hd__o21a_1
XFILLER_117_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15348_ _15348_/A vssd1 vssd1 vccd1 vccd1 _18723_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_25_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19612_/CLK sky130_fd_sc_hd__clkbuf_16
X_18067_ _19809_/Q _18067_/B _18067_/C vssd1 vssd1 vccd1 vccd1 _18069_/B sky130_fd_sc_hd__and3_1
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10050__A3 _10049_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15279_ _15279_/A vssd1 vssd1 vccd1 vccd1 _18693_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17018_ _17018_/A vssd1 vssd1 vccd1 vccd1 _19413_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10338__A1 _19061_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16898__S _16902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12504__B _12505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ _11148_/A _12497_/A vssd1 vssd1 vccd1 vccd1 _11147_/A sky130_fd_sc_hd__nand2_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10305__A _11166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09771_ _18610_/Q _19299_/Q _10010_/S vssd1 vssd1 vccd1 vccd1 _09771_/X sky130_fd_sc_hd__mux2_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ _19589_/CLK _18969_/D vssd1 vssd1 vccd1 vccd1 _18969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15307__S _15311_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14788__A0 _18433_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09205_ _09861_/A vssd1 vssd1 vccd1 vccd1 _09856_/A sky130_fd_sc_hd__buf_2
XANTENNA__15977__S _15983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11369__A3 _11593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09967__B1 _09892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09136_ _19692_/Q vssd1 vssd1 vccd1 vccd1 _10960_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10121__S0 _10011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10672__S1 _10616_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14712__B1 _14708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_8_0_clock clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_8_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_77_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09969_ _09969_/A _09969_/B vssd1 vssd1 vccd1 vccd1 _09969_/X sky130_fd_sc_hd__or2_1
XANTENNA__15217__S _15217_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11829__A1 _15262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ _12982_/B _12982_/C _12979_/Y vssd1 vssd1 vccd1 vccd1 _18307_/D sky130_fd_sc_hd__o21a_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10188__S0 _09721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _11984_/A _11984_/D vssd1 vssd1 vccd1 vccd1 _11957_/B sky130_fd_sc_hd__nand2_1
XFILLER_18_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11046__A _11046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _14553_/A _14648_/X _14649_/X input41/X vssd1 vssd1 vccd1 vccd1 _17775_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _12473_/A _12173_/A _12023_/B _11514_/A vssd1 vssd1 vccd1 vccd1 _11913_/A
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13601_ _13765_/S vssd1 vssd1 vccd1 vccd1 _13757_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_26_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10813_ _10813_/A _10813_/B vssd1 vssd1 vccd1 vccd1 _10813_/X sky130_fd_sc_hd__and2_1
XANTENNA__12254__A1 _13523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17717__A0 _12656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14581_ _18549_/Q _14577_/X _14580_/X _14573_/X vssd1 vssd1 vccd1 vccd1 _18549_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _12117_/B vssd1 vssd1 vccd1 vccd1 _12095_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_14_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09655__C1 _09708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16320_ _16342_/A vssd1 vssd1 vccd1 vccd1 _16329_/S sky130_fd_sc_hd__clkbuf_4
X_13532_ _13532_/A _13536_/A vssd1 vssd1 vccd1 vccd1 _13537_/A sky130_fd_sc_hd__nor2_2
XFILLER_159_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10744_ _18759_/Q _18988_/Q _18919_/Q _19217_/Q _10858_/A _10740_/X vssd1 vssd1 vccd1
+ vccd1 _10745_/B sky130_fd_sc_hd__mux4_1
XFILLER_159_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15887__S _15891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16251_ _16087_/X _19099_/Q _16257_/S vssd1 vssd1 vccd1 vccd1 _16252_/A sky130_fd_sc_hd__mux2_1
X_13463_ _13463_/A vssd1 vssd1 vccd1 vccd1 _18391_/D sky130_fd_sc_hd__clkbuf_1
X_10675_ _10875_/A _10675_/B vssd1 vssd1 vccd1 vccd1 _10675_/X sky130_fd_sc_hd__or2_1
X_15202_ _15202_/A vssd1 vssd1 vccd1 vccd1 _18670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12414_ _18379_/Q _12414_/B vssd1 vssd1 vccd1 vccd1 _12439_/B sky130_fd_sc_hd__and2_1
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16182_ _16182_/A vssd1 vssd1 vccd1 vccd1 _19064_/D sky130_fd_sc_hd__clkbuf_1
X_13394_ _19820_/Q vssd1 vssd1 vccd1 vccd1 _18102_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_138_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15133_ _16639_/A vssd1 vssd1 vccd1 vccd1 _15133_/X sky130_fd_sc_hd__buf_2
XFILLER_5_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12345_ _12345_/A vssd1 vssd1 vccd1 vccd1 _12345_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09973__A3 _09972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13506__A1 _13399_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09186__A _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15064_ _11542_/X _15062_/X _15063_/X vssd1 vssd1 vccd1 vccd1 _16737_/A sky130_fd_sc_hd__o21a_4
X_12276_ _19751_/Q _12116_/X _12271_/X _12275_/Y vssd1 vssd1 vccd1 vccd1 _17900_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_5_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09805__S0 _09803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14015_ _18433_/Q _14014_/X _14032_/S vssd1 vssd1 vccd1 vccd1 _14016_/A sky130_fd_sc_hd__mux2_1
X_11227_ _11227_/A _11229_/A _11227_/C vssd1 vssd1 vccd1 vccd1 _11227_/Y sky130_fd_sc_hd__nand3_1
X_19872_ _19872_/CLK _19872_/D vssd1 vssd1 vccd1 vccd1 _19872_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10125__A _10125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10415__S1 _09142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12190__A0 _12185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14820__A _16670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09914__A _09914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18823_ _19539_/CLK _18823_/D vssd1 vssd1 vccd1 vccd1 _18823_/Q sky130_fd_sc_hd__dfxtp_1
X_11158_ _09172_/A _11157_/X _09184_/A vssd1 vssd1 vccd1 vccd1 _11158_/X sky130_fd_sc_hd__a21o_1
XFILLER_95_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10109_ _19616_/Q _19454_/Q _18900_/Q _18670_/Q _10154_/S _10103_/A vssd1 vssd1 vccd1
+ vccd1 _10110_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12340__A _18376_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18754_ _19597_/CLK _18754_/D vssd1 vssd1 vccd1 vccd1 _18754_/Q sky130_fd_sc_hd__dfxtp_1
X_15966_ _14729_/X _18983_/Q _15972_/S vssd1 vssd1 vccd1 vccd1 _15967_/A sky130_fd_sc_hd__mux2_1
X_11089_ _09170_/A _11088_/X _09454_/A vssd1 vssd1 vccd1 vccd1 _11089_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17705_ _19677_/Q _17704_/X _17718_/S vssd1 vssd1 vccd1 vccd1 _17706_/A sky130_fd_sc_hd__mux2_1
X_14917_ _16696_/A vssd1 vssd1 vccd1 vccd1 _16800_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18685_ _19472_/CLK _18685_/D vssd1 vssd1 vccd1 vccd1 _18685_/Q sky130_fd_sc_hd__dfxtp_1
X_15897_ _15897_/A vssd1 vssd1 vccd1 vccd1 _18951_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17636_ _13212_/X _17634_/Y _17658_/S vssd1 vssd1 vccd1 vccd1 _17636_/X sky130_fd_sc_hd__mux2_1
X_14848_ _14847_/X _18597_/Q _14880_/S vssd1 vssd1 vccd1 vccd1 _14849_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15431__A1 _15159_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17567_ _17567_/A vssd1 vssd1 vccd1 vccd1 _19642_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09646__C1 _09689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14779_ _14776_/X _14777_/X _14893_/A vssd1 vssd1 vccd1 vccd1 _14779_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13171__A _13171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19306_ _19628_/CLK _19306_/D vssd1 vssd1 vccd1 vccd1 _19306_/Q sky130_fd_sc_hd__dfxtp_1
X_16518_ _16518_/A vssd1 vssd1 vccd1 vccd1 _19216_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17184__A1 _13279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17498_ _17520_/A vssd1 vssd1 vccd1 vccd1 _17507_/S sky130_fd_sc_hd__buf_2
XFILLER_31_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19237_ _19722_/CLK _19237_/D vssd1 vssd1 vccd1 vccd1 _19237_/Q sky130_fd_sc_hd__dfxtp_1
X_16449_ _16058_/X _19186_/Q _16453_/S vssd1 vssd1 vccd1 vccd1 _16450_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19168_ _19618_/CLK _19168_/D vssd1 vssd1 vccd1 vccd1 _19168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18119_ _19827_/Q _18119_/B _18119_/C vssd1 vssd1 vccd1 vccd1 _18120_/C sky130_fd_sc_hd__and3_1
XFILLER_118_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19099_ _19612_/CLK _19099_/D vssd1 vssd1 vccd1 vccd1 _19099_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10654__S1 _09353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15498__A1 _15497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10406__S1 _09602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09823_ _09865_/A vssd1 vssd1 vccd1 vccd1 _09952_/S sky130_fd_sc_hd__buf_2
XFILLER_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10192__C1 _09395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10731__B2 _18433_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09754_ _11222_/A _12500_/A vssd1 vssd1 vccd1 vccd1 _09756_/B sky130_fd_sc_hd__or2_1
XFILLER_55_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13681__A0 _12262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09685_ _09402_/A _09669_/X _09684_/X vssd1 vssd1 vccd1 vccd1 _09685_/X sky130_fd_sc_hd__a21o_2
XFILLER_104_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17252__S _17258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10590__S0 _10511_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10460_ _10461_/A _12480_/A vssd1 vssd1 vccd1 vccd1 _10462_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11724__A1_N _11820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09119_ _09119_/A _09119_/B vssd1 vssd1 vccd1 vccd1 _13578_/A sky130_fd_sc_hd__nand2_8
XFILLER_109_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10391_ _10239_/X _10388_/Y _10390_/Y _10496_/A vssd1 vssd1 vccd1 vccd1 _10391_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12130_ _14155_/A _14168_/A vssd1 vssd1 vccd1 vccd1 _12131_/D sky130_fd_sc_hd__or2_1
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12144__B _19746_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10970__A1 _09169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17427__S _17435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12061_ _11135_/A _18505_/Q _12177_/A vssd1 vssd1 vccd1 vccd1 _13603_/A sky130_fd_sc_hd__mux2_4
XANTENNA__15736__A _17391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11012_ _18981_/Q _11012_/B _11012_/C vssd1 vssd1 vccd1 vccd1 _11012_/X sky130_fd_sc_hd__or3_1
XFILLER_77_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15820_ _15820_/A vssd1 vssd1 vccd1 vccd1 _18917_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _15751_/A vssd1 vssd1 vccd1 vccd1 _18886_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12963_ _18298_/Q _12961_/A _12962_/X vssd1 vssd1 vccd1 vccd1 _18298_/D sky130_fd_sc_hd__o21ba_1
XANTENNA__13672__A0 _12424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14702_ _14802_/A _14701_/Y _19080_/Q _11381_/C vssd1 vssd1 vccd1 vccd1 _14703_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_166_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ _11866_/B _11913_/Y _11970_/A vssd1 vssd1 vccd1 vccd1 _11915_/B sky130_fd_sc_hd__a21o_1
X_18470_ _19080_/CLK _18470_/D vssd1 vssd1 vccd1 vccd1 _18470_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11683__C1 _11997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15682_ _18856_/Q _15513_/X _15686_/S vssd1 vssd1 vccd1 vccd1 _15683_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12894_ _12904_/A _12894_/B _12894_/C vssd1 vssd1 vccd1 vccd1 _18277_/D sky130_fd_sc_hd__nor3_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _17421_/A vssd1 vssd1 vccd1 vccd1 _19577_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _14648_/A vssd1 vssd1 vccd1 vccd1 _14633_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12227__A1 _14568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _11810_/A _13984_/B _11844_/X vssd1 vssd1 vccd1 vccd1 _11846_/B sky130_fd_sc_hd__a21oi_2
XFILLER_33_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output104_A _11899_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _16790_/X _19547_/Q _17352_/S vssd1 vssd1 vccd1 vccd1 _17353_/A sky130_fd_sc_hd__mux2_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14572_/B vssd1 vssd1 vccd1 vccd1 _14564_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _11776_/A vssd1 vssd1 vccd1 vccd1 _11970_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16303_ _16058_/X _19122_/Q _16307_/S vssd1 vssd1 vccd1 vccd1 _16304_/A sky130_fd_sc_hd__mux2_1
X_13515_ _14589_/B vssd1 vssd1 vccd1 vccd1 _14526_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10727_ _19410_/Q _19186_/Q _19703_/Q _19154_/Q _10724_/X _10726_/X vssd1 vssd1 vccd1
+ vccd1 _10727_/X sky130_fd_sc_hd__mux4_1
X_17283_ _19516_/Q _16689_/X _17291_/S vssd1 vssd1 vccd1 vccd1 _17284_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11450__A2 _13108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14495_ _14495_/A vssd1 vssd1 vccd1 vccd1 _18517_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16506__S _16514_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19022_ _19638_/CLK _19022_/D vssd1 vssd1 vccd1 vccd1 _19022_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15410__S _15410_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16234_ _16234_/A vssd1 vssd1 vccd1 vccd1 _19091_/D sky130_fd_sc_hd__clkbuf_1
X_13446_ _13446_/A vssd1 vssd1 vccd1 vccd1 _18383_/D sky130_fd_sc_hd__clkbuf_1
X_10658_ _10589_/A _10643_/X _10657_/X vssd1 vssd1 vccd1 vccd1 _10658_/X sky130_fd_sc_hd__a21o_2
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16165_ _16165_/A vssd1 vssd1 vccd1 vccd1 _19056_/D sky130_fd_sc_hd__clkbuf_1
X_13377_ _18376_/Q _13413_/B vssd1 vssd1 vccd1 vccd1 _13377_/X sky130_fd_sc_hd__or2_1
XANTENNA__09628__B _12503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09800__C1 _09249_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12335__A _19753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10589_ _10589_/A _10589_/B _10589_/C vssd1 vssd1 vccd1 vccd1 _10589_/X sky130_fd_sc_hd__or3_2
XFILLER_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15116_ _15116_/A vssd1 vssd1 vccd1 vccd1 _15116_/X sky130_fd_sc_hd__buf_2
XFILLER_127_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12328_ _12328_/A vssd1 vssd1 vccd1 vccd1 _12423_/S sky130_fd_sc_hd__clkbuf_4
X_16096_ _16806_/A vssd1 vssd1 vccd1 vccd1 _16096_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15047_ input22/X _14960_/A _15000_/X vssd1 vssd1 vccd1 vccd1 _15047_/X sky130_fd_sc_hd__a21o_1
X_12259_ _18513_/Q _12259_/B _12259_/C vssd1 vssd1 vccd1 vccd1 _12259_/X sky130_fd_sc_hd__or3_1
XFILLER_68_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19855_ _19855_/CLK _19855_/D vssd1 vssd1 vccd1 vccd1 _19855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11061__S1 _09480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18806_ _19003_/CLK _18806_/D vssd1 vssd1 vccd1 vccd1 _18806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19786_ _19786_/CLK _19786_/D vssd1 vssd1 vccd1 vccd1 _19786_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_23_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16998_ _16998_/A vssd1 vssd1 vccd1 vccd1 _19404_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18737_ _19452_/CLK _18737_/D vssd1 vssd1 vccd1 vccd1 _18737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15949_ _15949_/A vssd1 vssd1 vccd1 vccd1 _18975_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16477__A _16488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09470_ _09434_/X _09463_/X _09465_/X _09469_/X _09246_/A vssd1 vssd1 vccd1 vccd1
+ _09470_/X sky130_fd_sc_hd__a311o_2
XFILLER_92_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18668_ _19642_/CLK _18668_/D vssd1 vssd1 vccd1 vccd1 _18668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17619_ _19662_/Q _17618_/X _17625_/S vssd1 vssd1 vccd1 vccd1 _17620_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_178_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18599_ _19513_/CLK _18599_/D vssd1 vssd1 vccd1 vccd1 _18599_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17157__A1 _13197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16416__S _16424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15320__S _15322_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09819__A _09819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12245__A _12246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09554__A _09554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09806_ _09819_/A _09806_/B vssd1 vssd1 vccd1 vccd1 _09806_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13103__C1 _13102_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12457__A1 _19759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ _18779_/Q _19008_/Q _18939_/Q _19237_/Q _09734_/X _10186_/A vssd1 vssd1 vccd1
+ vccd1 _09737_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15291__A _15337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09668_ _09661_/A _09667_/X _09412_/A vssd1 vssd1 vccd1 vccd1 _09668_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_27_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13523__B _13523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10483__A3 _10482_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ _10279_/S vssd1 vssd1 vccd1 vccd1 _09600_/A sky130_fd_sc_hd__buf_2
XFILLER_43_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _12715_/B _11979_/A _12219_/S _11624_/Y vssd1 vssd1 vccd1 vccd1 _11630_/X
+ sky130_fd_sc_hd__or4b_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11968__A0 _12480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11561_ _11561_/A vssd1 vssd1 vccd1 vccd1 _12017_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14635__A _14654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13300_ _18318_/Q _13178_/A _12664_/A _19807_/Q _13299_/X vssd1 vssd1 vccd1 vccd1
+ _13300_/X sky130_fd_sc_hd__a221o_1
XFILLER_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15230__S _15233_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10512_ _10245_/A _10511_/X _10593_/A vssd1 vssd1 vccd1 vccd1 _10512_/X sky130_fd_sc_hd__a21o_1
X_14280_ _13823_/A _13949_/B _14279_/X _14115_/X vssd1 vssd1 vccd1 vccd1 _14280_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_156_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11492_ _14589_/A _14587_/A vssd1 vssd1 vccd1 vccd1 _13524_/C sky130_fd_sc_hd__or2_2
XFILLER_137_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13231_ _18358_/Q _13246_/B vssd1 vssd1 vccd1 vccd1 _13231_/X sky130_fd_sc_hd__or2_1
XFILLER_137_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10443_ _19641_/Q _19058_/Q _19095_/Q _18701_/Q _09673_/S _09486_/X vssd1 vssd1 vccd1
+ vccd1 _10443_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11196__A1 _09403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09484__S1 _09483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13162_ _19794_/Q _12518_/X _12522_/X _18305_/Q _13161_/X vssd1 vssd1 vccd1 vccd1
+ _13163_/B sky130_fd_sc_hd__a221o_2
XANTENNA_input65_A io_ibus_inst[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ _19515_/Q _19129_/Q _19579_/Q _18735_/Q _09448_/S _10349_/A vssd1 vssd1 vccd1
+ vccd1 _10375_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10943__A1 _10950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14134__A1 _18440_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12113_ _12089_/A _12089_/B _12086_/A vssd1 vssd1 vccd1 vccd1 _12114_/B sky130_fd_sc_hd__a21o_1
XFILLER_152_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13093_ _13093_/A vssd1 vssd1 vccd1 vccd1 _18342_/D sky130_fd_sc_hd__clkbuf_1
X_17970_ _19774_/Q _17971_/C _19775_/Q vssd1 vssd1 vccd1 vccd1 _17972_/B sky130_fd_sc_hd__a21oi_1
XFILLER_152_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12044_ _12067_/B _12044_/B vssd1 vssd1 vccd1 vccd1 _12044_/X sky130_fd_sc_hd__xor2_1
X_16921_ _16977_/A vssd1 vssd1 vccd1 vccd1 _16990_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_104_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17084__A0 _16771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19640_ _19640_/CLK _19640_/D vssd1 vssd1 vccd1 vccd1 _19640_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_5_0_clock clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
X_16852_ _19340_/Q _16645_/X _16858_/S vssd1 vssd1 vccd1 vccd1 _16853_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15803_ _15803_/A vssd1 vssd1 vccd1 vccd1 _18910_/D sky130_fd_sc_hd__clkbuf_1
X_16783_ _16783_/A vssd1 vssd1 vccd1 vccd1 _19318_/D sky130_fd_sc_hd__clkbuf_1
X_19571_ _19571_/CLK _19571_/D vssd1 vssd1 vccd1 vccd1 _19571_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12448__A1 _14324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13995_ _13992_/Y _13994_/Y _13995_/S vssd1 vssd1 vccd1 vccd1 _13995_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15734_ _18880_/Q _15589_/X _15734_/S vssd1 vssd1 vccd1 vccd1 _15735_/A sky130_fd_sc_hd__mux2_1
X_18522_ _18564_/CLK _18522_/D vssd1 vssd1 vccd1 vccd1 _18522_/Q sky130_fd_sc_hd__dfxtp_1
X_12946_ _18292_/Q _18291_/Q _12946_/C vssd1 vssd1 vccd1 vccd1 _12952_/C sky130_fd_sc_hd__and3_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09864__A2 _09854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15665_ _15721_/A vssd1 vssd1 vccd1 vccd1 _15734_/S sky130_fd_sc_hd__buf_8
XFILLER_34_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18453_ _19468_/CLK _18453_/D vssd1 vssd1 vccd1 vccd1 _18453_/Q sky130_fd_sc_hd__dfxtp_4
X_12877_ _12897_/A _12883_/C vssd1 vssd1 vccd1 vccd1 _12877_/Y sky130_fd_sc_hd__nor2_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _14616_/A vssd1 vssd1 vccd1 vccd1 _18559_/D sky130_fd_sc_hd__clkbuf_1
X_17404_ _17461_/S vssd1 vssd1 vccd1 vccd1 _17413_/S sky130_fd_sc_hd__buf_2
X_18384_ _19472_/CLK _18384_/D vssd1 vssd1 vccd1 vccd1 _18384_/Q sky130_fd_sc_hd__dfxtp_1
X_11828_ _11888_/C _11825_/X _11826_/Y _11827_/X vssd1 vssd1 vccd1 vccd1 _11828_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15596_ _15596_/A vssd1 vssd1 vccd1 vccd1 _18817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16744__B _17064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _16765_/X _19539_/Q _17341_/S vssd1 vssd1 vccd1 vccd1 _17336_/A sky130_fd_sc_hd__mux2_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _14547_/A _14551_/B vssd1 vssd1 vccd1 vccd1 _14547_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11759_ _18353_/Q _11759_/B vssd1 vssd1 vccd1 vccd1 _11759_/X sky130_fd_sc_hd__and2_1
XFILLER_53_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17266_ _17266_/A vssd1 vssd1 vccd1 vccd1 _19508_/D sky130_fd_sc_hd__clkbuf_1
X_14478_ _14591_/B vssd1 vssd1 vccd1 vccd1 _14487_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_146_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19005_ _19395_/CLK _19005_/D vssd1 vssd1 vccd1 vccd1 _19005_/Q sky130_fd_sc_hd__dfxtp_1
X_16217_ _16217_/A vssd1 vssd1 vccd1 vccd1 _19083_/D sky130_fd_sc_hd__clkbuf_1
X_13429_ _19500_/Q _13418_/S _12671_/A _18688_/Q vssd1 vssd1 vccd1 vccd1 _13429_/X
+ sky130_fd_sc_hd__a22o_1
X_17197_ _17197_/A vssd1 vssd1 vccd1 vccd1 _19485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16148_ _16045_/X _19049_/Q _16150_/S vssd1 vssd1 vccd1 vccd1 _16149_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17067__S _17075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16079_ _16079_/A vssd1 vssd1 vccd1 vccd1 _19027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12687__A1 _13112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15095__B _15095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10147__C1 _09404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17075__A0 _16758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10698__B1 _09407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19838_ _19838_/CLK _19838_/D vssd1 vssd1 vccd1 vccd1 _19838_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__10313__A _10313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13636__A0 _13658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 io_dbus_rdata[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
X_19769_ _19779_/CLK _19769_/D vssd1 vssd1 vccd1 vccd1 _19769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13100__A2 _12731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ _09522_/A vssd1 vssd1 vccd1 vccd1 _11110_/S sky130_fd_sc_hd__clkbuf_4
X_09453_ _09695_/A _09448_/X _09452_/X vssd1 vssd1 vccd1 vccd1 _09453_/X sky130_fd_sc_hd__a21o_1
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11144__A _12495_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09384_ _10068_/A vssd1 vssd1 vccd1 vccd1 _09385_/A sky130_fd_sc_hd__buf_2
XFILLER_40_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16146__S _16150_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09268__B _18533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16670__A _16670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09466__S1 _09142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12703__A _12703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10090_ _19649_/Q _19066_/Q _19103_/Q _18709_/Q _10153_/S _09769_/A vssd1 vssd1 vccd1
+ vccd1 _10090_/X sky130_fd_sc_hd__mux4_1
XFILLER_160_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10138__C1 _09395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11025__S1 _10920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13875__B1 _18428_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12800_ _12813_/D vssd1 vssd1 vccd1 vccd1 _18250_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13534__A _13542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13780_ _13770_/X _13777_/X _14121_/S vssd1 vssd1 vccd1 vccd1 _13780_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10992_ _10992_/A _10992_/B vssd1 vssd1 vccd1 vccd1 _10992_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12346__A1_N _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12731_ _12731_/A vssd1 vssd1 vccd1 vccd1 _12731_/X sky130_fd_sc_hd__buf_2
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10310__C1 _09562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17440__S _17446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15450_ _15472_/A vssd1 vssd1 vccd1 vccd1 _15459_/S sky130_fd_sc_hd__clkbuf_4
X_12662_ _13130_/A vssd1 vssd1 vccd1 vccd1 _13178_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14052__A0 _18435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _18479_/Q _18511_/Q _14410_/S vssd1 vssd1 vccd1 vccd1 _14402_/A sky130_fd_sc_hd__mux2_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11692_/A _11692_/B _11613_/C vssd1 vssd1 vccd1 vccd1 _11613_/X sky130_fd_sc_hd__or3_1
XFILLER_30_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15381_ _15381_/A vssd1 vssd1 vccd1 vccd1 _18738_/D sky130_fd_sc_hd__clkbuf_1
X_12593_ _19809_/Q _12518_/X _12522_/X _18320_/Q _12592_/X vssd1 vssd1 vccd1 vccd1
+ _12594_/B sky130_fd_sc_hd__a221o_2
XANTENNA__16056__S _16065_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17120_ _17120_/A vssd1 vssd1 vccd1 vccd1 _19459_/D sky130_fd_sc_hd__clkbuf_1
X_14332_ _14332_/A _14332_/B vssd1 vssd1 vccd1 vccd1 _14332_/X sky130_fd_sc_hd__or2_1
X_11544_ _11542_/X _13578_/A _14032_/S vssd1 vssd1 vccd1 vccd1 _11545_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17051_ _17051_/A vssd1 vssd1 vccd1 vccd1 _19428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14263_ _11602_/Y _14265_/A _14088_/A _14262_/X vssd1 vssd1 vccd1 vccd1 _14263_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11475_ _11475_/A _11585_/B _11642_/C vssd1 vssd1 vccd1 vccd1 _13583_/B sky130_fd_sc_hd__or3_2
XFILLER_125_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16002_ _16002_/A vssd1 vssd1 vccd1 vccd1 _18999_/D sky130_fd_sc_hd__clkbuf_1
X_13214_ _13185_/X _13212_/X _13213_/X _13167_/X vssd1 vssd1 vccd1 vccd1 _18356_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_137_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10426_ _09689_/A _10416_/X _10420_/X _10425_/X _09133_/A vssd1 vssd1 vccd1 vccd1
+ _10426_/X sky130_fd_sc_hd__a311o_4
XFILLER_100_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14194_ _14182_/A _14191_/X _14193_/Y _13950_/A vssd1 vssd1 vccd1 vccd1 _14194_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10916__A1 _10956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_126_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ _19857_/Q _12604_/A _12583_/A _19825_/Q vssd1 vssd1 vccd1 vccd1 _13145_/X
+ sky130_fd_sc_hd__a22o_1
X_10357_ _10928_/A vssd1 vssd1 vccd1 vccd1 _10866_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13315__C1 _13282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _17954_/B _17954_/C _19769_/Q vssd1 vssd1 vccd1 vccd1 _17955_/B sky130_fd_sc_hd__a21oi_1
X_13076_ _13324_/A _18626_/Q vssd1 vssd1 vccd1 vccd1 _13076_/Y sky130_fd_sc_hd__nand2_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _10288_/A _10288_/B vssd1 vssd1 vccd1 vccd1 _10288_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16904_ _16904_/A vssd1 vssd1 vccd1 vccd1 _16913_/S sky130_fd_sc_hd__buf_6
X_12027_ _11474_/A _12026_/X _12126_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _12028_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_17884_ _17890_/A _17884_/B vssd1 vssd1 vccd1 vccd1 _17885_/A sky130_fd_sc_hd__and2_1
XFILLER_39_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19623_ _19722_/CLK _19623_/D vssd1 vssd1 vccd1 vccd1 _19623_/Q sky130_fd_sc_hd__dfxtp_1
X_16835_ _16835_/A vssd1 vssd1 vccd1 vccd1 _16835_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19554_ _19554_/CLK _19554_/D vssd1 vssd1 vccd1 vccd1 _19554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16766_ _16765_/X _19313_/Q _16775_/S vssd1 vssd1 vccd1 vccd1 _16767_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13978_ _14262_/A vssd1 vssd1 vccd1 vccd1 _13978_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14830__A2 _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18505_ _18506_/CLK _18505_/D vssd1 vssd1 vccd1 vccd1 _18505_/Q sky130_fd_sc_hd__dfxtp_1
X_12929_ _12897_/B _12933_/D _18287_/Q vssd1 vssd1 vccd1 vccd1 _12931_/B sky130_fd_sc_hd__a21oi_1
X_15717_ _18872_/Q _15564_/X _15719_/S vssd1 vssd1 vccd1 vccd1 _15718_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13163__B _13163_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19485_ _19488_/CLK _19485_/D vssd1 vssd1 vccd1 vccd1 _19485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16697_ _19292_/Q _16696_/X _16703_/S vssd1 vssd1 vccd1 vccd1 _16698_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10279__S _10279_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17350__S _17352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18436_ _18818_/CLK _18436_/D vssd1 vssd1 vccd1 vccd1 _18436_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_62_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15648_ _15648_/A vssd1 vssd1 vccd1 vccd1 _18841_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18367_ _18402_/CLK _18367_/D vssd1 vssd1 vccd1 vccd1 _18367_/Q sky130_fd_sc_hd__dfxtp_1
X_15579_ _15579_/A vssd1 vssd1 vccd1 vccd1 _18812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17318_ _17318_/A vssd1 vssd1 vccd1 vccd1 _19532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18298_ _18298_/CLK _18298_/D vssd1 vssd1 vccd1 vccd1 _18298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17249_ _17317_/S vssd1 vssd1 vccd1 vccd1 _17258_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12109__A0 _11137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10383__A2 _10373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11139__A _11139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17525__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09620__S1 _11189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09832__A _10068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13609__A0 _14126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15045__S _15056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14282__A0 _18452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09505_ _18783_/Q _19012_/Q _18943_/Q _19241_/Q _10277_/S _09501_/A vssd1 vssd1 vccd1
+ vccd1 _09506_/B sky130_fd_sc_hd__mux4_1
XFILLER_112_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11191__S0 _10185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _10905_/S vssd1 vssd1 vccd1 vccd1 _10982_/S sky130_fd_sc_hd__clkbuf_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _18880_/Q _19338_/Q _09367_/S vssd1 vssd1 vccd1 vccd1 _09368_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09298_ _18578_/Q vssd1 vssd1 vccd1 vccd1 _14572_/A sky130_fd_sc_hd__inv_2
XFILLER_138_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11260_ _11244_/A _10601_/X _11080_/B _11080_/C vssd1 vssd1 vccd1 vccd1 _11260_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10211_ _19518_/Q _19132_/Q _19582_/Q _18738_/Q _10094_/A _09978_/A vssd1 vssd1 vccd1
+ vccd1 _10212_/B sky130_fd_sc_hd__mux4_1
XFILLER_134_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13529__A _13529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12433__A _19758_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11191_ _18781_/Q _19010_/Q _18941_/Q _19239_/Q _10185_/S _09728_/A vssd1 vssd1 vccd1
+ vccd1 _11191_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10142_ _10144_/A _10141_/X _09414_/A vssd1 vssd1 vccd1 vccd1 _10142_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13248__B _18629_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17435__S _17435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10073_ _19263_/Q _19034_/Q _18965_/Q _19359_/Q _10114_/S _09984_/A vssd1 vssd1 vccd1
+ vccd1 _10074_/B sky130_fd_sc_hd__mux4_1
X_14950_ _16705_/A vssd1 vssd1 vccd1 vccd1 _16809_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09611__S1 _09610_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13901_ _14130_/A _13901_/B vssd1 vssd1 vccd1 vccd1 _13908_/B sky130_fd_sc_hd__nor2_1
X_14881_ _14881_/A vssd1 vssd1 vccd1 vccd1 _18600_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input28_A io_dbus_rdata[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16620_ _16620_/A vssd1 vssd1 vccd1 vccd1 _19265_/D sky130_fd_sc_hd__clkbuf_1
X_13832_ _13832_/A vssd1 vssd1 vccd1 vccd1 _14328_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16551_ _16551_/A vssd1 vssd1 vccd1 vccd1 _19231_/D sky130_fd_sc_hd__clkbuf_1
X_13763_ _13753_/X _13760_/X _13918_/S vssd1 vssd1 vccd1 vccd1 _13763_/X sky130_fd_sc_hd__a21o_1
X_10975_ _10992_/A _10975_/B vssd1 vssd1 vccd1 vccd1 _10975_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ _13108_/B _12714_/B _13108_/A vssd1 vssd1 vccd1 vccd1 _12714_/X sky130_fd_sc_hd__or3b_1
X_15502_ _15502_/A vssd1 vssd1 vccd1 vccd1 _18788_/D sky130_fd_sc_hd__clkbuf_1
X_16482_ _16106_/X _19201_/Q _16486_/S vssd1 vssd1 vccd1 vccd1 _16483_/A sky130_fd_sc_hd__mux2_1
X_19270_ _19579_/CLK _19270_/D vssd1 vssd1 vccd1 vccd1 _19270_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_52_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13694_ _14036_/S vssd1 vssd1 vccd1 vccd1 _14019_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18221_ _18221_/A _18221_/B vssd1 vssd1 vccd1 vccd1 _19861_/D sky130_fd_sc_hd__nor2_1
X_15433_ _18760_/Q _15162_/X _15437_/S vssd1 vssd1 vccd1 vccd1 _15434_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12645_ _19679_/Q _12624_/A _12674_/A _18403_/Q vssd1 vssd1 vccd1 vccd1 _12645_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13711__B _13711_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09678__S1 _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18152_ _19837_/Q _18150_/B _18151_/Y vssd1 vssd1 vccd1 vccd1 _19837_/D sky130_fd_sc_hd__o21a_1
X_15364_ _15410_/S vssd1 vssd1 vccd1 vccd1 _15373_/S sky130_fd_sc_hd__buf_4
X_12576_ _12600_/A vssd1 vssd1 vccd1 vccd1 _13297_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09452__B1 _09454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10598__C1 _09392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10062__A1 _09892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14315_ _13949_/A _13851_/X _14314_/Y _14054_/A vssd1 vssd1 vccd1 vccd1 _14315_/X
+ sky130_fd_sc_hd__o211a_1
X_17103_ _17103_/A vssd1 vssd1 vccd1 vccd1 _19451_/D sky130_fd_sc_hd__clkbuf_1
X_18083_ _18086_/B _18086_/C _18082_/X vssd1 vssd1 vccd1 vccd1 _18083_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11527_ _11599_/A vssd1 vssd1 vccd1 vccd1 _12505_/B sky130_fd_sc_hd__buf_2
X_15295_ _15295_/A vssd1 vssd1 vccd1 vccd1 _18700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16514__S _16514_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10128__A _10328_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17034_ _19421_/Q _16699_/X _17036_/S vssd1 vssd1 vccd1 vccd1 _17035_/A sky130_fd_sc_hd__mux2_1
X_14246_ _12265_/Y _14102_/X _14245_/X vssd1 vssd1 vccd1 vccd1 _14246_/X sky130_fd_sc_hd__a21bo_1
X_11458_ _11458_/A vssd1 vssd1 vccd1 vccd1 _15093_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10409_ _10398_/X _10408_/X _10494_/A vssd1 vssd1 vccd1 vccd1 _10409_/X sky130_fd_sc_hd__mux2_4
X_14177_ _13977_/A _14176_/B _14040_/A vssd1 vssd1 vccd1 vccd1 _14177_/X sky130_fd_sc_hd__o21a_1
X_11389_ _11388_/Y _18421_/Q _14900_/B vssd1 vssd1 vccd1 vccd1 _14801_/A sky130_fd_sc_hd__mux2_4
XFILLER_124_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _12863_/B _13126_/X _13127_/X _18350_/Q vssd1 vssd1 vccd1 vccd1 _13128_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ _19597_/CLK _18985_/D vssd1 vssd1 vccd1 vccd1 _18985_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12062__B _13603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14500__A1 _19758_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17936_ _19764_/Q _19763_/Q _19762_/Q _17936_/D vssd1 vssd1 vccd1 vccd1 _17946_/D
+ sky130_fd_sc_hd__and4_1
X_13059_ _13069_/D vssd1 vssd1 vccd1 vccd1 _13067_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17867_ _17867_/A vssd1 vssd1 vccd1 vccd1 _19734_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_2_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_19606_ _19659_/CLK _19606_/D vssd1 vssd1 vccd1 vccd1 _19606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16818_ _16818_/A vssd1 vssd1 vccd1 vccd1 _19329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17798_ _17798_/A vssd1 vssd1 vccd1 vccd1 _19701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19537_ _19537_/CLK _19537_/D vssd1 vssd1 vccd1 vccd1 _19537_/Q sky130_fd_sc_hd__dfxtp_1
X_16749_ _16749_/A vssd1 vssd1 vccd1 vccd1 _16749_/X sky130_fd_sc_hd__buf_2
XANTENNA__11617__A2 _11940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17202__A0 _19487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19468_ _19468_/CLK _19468_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09221_ _09856_/A _09221_/B vssd1 vssd1 vccd1 vccd1 _09221_/X sky130_fd_sc_hd__or2_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18419_ _18509_/CLK _18419_/D vssd1 vssd1 vccd1 vccd1 _18419_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_50_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19399_ _19657_/CLK _19399_/D vssd1 vssd1 vccd1 vccd1 _19399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09152_ _09152_/A vssd1 vssd1 vccd1 vccd1 _10605_/S sky130_fd_sc_hd__buf_2
XFILLER_148_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09083_ _18560_/Q vssd1 vssd1 vccd1 vccd1 _11320_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16424__S _16424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18205__A _18205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput70 io_irq_spi_irq vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11553__A1 _11552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10987__S0 _10905_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09985_ _18775_/Q _19004_/Q _18935_/Q _19233_/Q _09983_/X _09984_/X vssd1 vssd1 vccd1
+ vccd1 _09986_/B sky130_fd_sc_hd__mux4_1
XFILLER_130_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15564__A _16819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09562__A _09708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10760_ _10850_/A _10760_/B vssd1 vssd1 vccd1 vccd1 _10760_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09682__B1 _09681_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10911__S0 _10909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09419_ _09814_/A _09419_/B vssd1 vssd1 vccd1 vccd1 _09419_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_4_0_clock clkbuf_4_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_4_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10691_ _09273_/A _10681_/X _10690_/X _09280_/A _18433_/Q vssd1 vssd1 vccd1 vccd1
+ _10691_/X sky130_fd_sc_hd__a32o_2
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12430_ _12430_/A _12430_/B vssd1 vssd1 vccd1 vccd1 _12431_/B sky130_fd_sc_hd__nand2_2
XFILLER_139_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13230__B2 _18627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12361_ _12361_/A _12387_/C vssd1 vssd1 vccd1 vccd1 _12386_/B sky130_fd_sc_hd__and2_1
XFILLER_148_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16334__S _16340_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14643__A _18205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14100_ _11978_/X _14070_/X _14098_/X _14099_/X vssd1 vssd1 vccd1 vccd1 _14100_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__13518__C1 _13542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_6_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19546_/CLK sky130_fd_sc_hd__clkbuf_16
X_11312_ _11501_/B _09119_/A _09119_/B vssd1 vssd1 vccd1 vccd1 _11580_/C sky130_fd_sc_hd__o21ai_1
X_15080_ _11497_/A _11591_/Y _15092_/S vssd1 vssd1 vccd1 vccd1 _15080_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12292_ _19752_/Q _12292_/B vssd1 vssd1 vccd1 vccd1 _12335_/C sky130_fd_sc_hd__and2_1
XFILLER_119_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14031_ _11880_/A _13933_/A _14030_/X vssd1 vssd1 vccd1 vccd1 _14031_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__17954__A _19769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11243_ _11242_/B _11242_/C _11242_/A vssd1 vssd1 vccd1 vccd1 _11243_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11544__A1 _13578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11174_ _09277_/A _11164_/X _11173_/X _09284_/A _18454_/Q vssd1 vssd1 vccd1 vccd1
+ _11199_/A sky130_fd_sc_hd__a32o_4
XANTENNA__14789__S _14893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17680__A0 _13294_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ _10125_/A vssd1 vssd1 vccd1 vccd1 _10125_/X sky130_fd_sc_hd__buf_2
XFILLER_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18770_ _19642_/CLK _18770_/D vssd1 vssd1 vccd1 vccd1 _18770_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14494__A0 _18517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15982_ _15982_/A vssd1 vssd1 vccd1 vccd1 _18990_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17721_ _17716_/A _17720_/C _18479_/Q vssd1 vssd1 vccd1 vccd1 _17721_/Y sky130_fd_sc_hd__o21ai_1
X_10056_ _09880_/A _10055_/X _10068_/A vssd1 vssd1 vccd1 vccd1 _10056_/X sky130_fd_sc_hd__a21o_1
X_14933_ _17701_/B _14932_/C _18477_/Q vssd1 vssd1 vccd1 vccd1 _14934_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__10504__C1 _09681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17652_ _13245_/X _17651_/Y _17658_/S vssd1 vssd1 vccd1 vccd1 _17652_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14864_ input5/X _14801_/A _14804_/A vssd1 vssd1 vccd1 vccd1 _14864_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10411__A _10412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16603_ _19257_/Q vssd1 vssd1 vccd1 vccd1 _16604_/A sky130_fd_sc_hd__clkbuf_1
X_13815_ _14034_/S _13818_/B vssd1 vssd1 vccd1 vccd1 _13816_/A sky130_fd_sc_hd__nand2_1
X_17583_ _17583_/A vssd1 vssd1 vccd1 vccd1 _19649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14795_ _17645_/A _14796_/B _14875_/A vssd1 vssd1 vccd1 vccd1 _14795_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19322_ _19581_/CLK _19322_/D vssd1 vssd1 vccd1 vccd1 _19322_/Q sky130_fd_sc_hd__dfxtp_1
X_13746_ _13668_/X _13661_/X _13747_/S vssd1 vssd1 vccd1 vccd1 _13746_/X sky130_fd_sc_hd__mux2_1
X_16534_ _19224_/Q _15532_/X _16536_/S vssd1 vssd1 vccd1 vccd1 _16535_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10958_ _11026_/A _10958_/B vssd1 vssd1 vccd1 vccd1 _10958_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19253_ _19285_/CLK _19253_/D vssd1 vssd1 vccd1 vccd1 _19253_/Q sky130_fd_sc_hd__dfxtp_1
X_13677_ _13664_/X _13675_/X _13965_/S vssd1 vssd1 vccd1 vccd1 _13677_/X sky130_fd_sc_hd__mux2_1
X_16465_ _16465_/A vssd1 vssd1 vccd1 vccd1 _19193_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12338__A _19685_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10889_ _19405_/Q _19181_/Q _19698_/Q _19149_/Q _10711_/A _10785_/X vssd1 vssd1 vccd1
+ vccd1 _10889_/X sky130_fd_sc_hd__mux4_2
XFILLER_32_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18204_ _19855_/Q _18201_/B _18203_/Y vssd1 vssd1 vccd1 vccd1 _19855_/D sky130_fd_sc_hd__o21a_1
X_12628_ _12628_/A vssd1 vssd1 vccd1 vccd1 _12629_/S sky130_fd_sc_hd__clkbuf_2
X_15416_ _15472_/A vssd1 vssd1 vccd1 vccd1 _15485_/S sky130_fd_sc_hd__buf_6
XANTENNA__13221__A1 _19667_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19184_ _19634_/CLK _19184_/D vssd1 vssd1 vccd1 vccd1 _19184_/Q sky130_fd_sc_hd__dfxtp_1
X_16396_ _19163_/Q _15542_/X _16402_/S vssd1 vssd1 vccd1 vccd1 _16397_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17499__A0 _19612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18135_ _18159_/A _18140_/C vssd1 vssd1 vccd1 vccd1 _18135_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12792__A1_N _11822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15347_ _18723_/Q _15146_/X _15351_/S vssd1 vssd1 vccd1 vccd1 _15348_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09520__S0 _10389_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12559_ _12514_/Y _12554_/X _12556_/X _12558_/X _18635_/Q vssd1 vssd1 vccd1 vccd1
+ _12559_/X sky130_fd_sc_hd__a32o_4
XANTENNA__14553__A _14553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16244__S _16246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18025__A _18033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18066_ _18067_/B _18067_/C _18065_/Y vssd1 vssd1 vccd1 vccd1 _19808_/D sky130_fd_sc_hd__o21a_1
X_15278_ _18693_/Q _15152_/X _15278_/S vssd1 vssd1 vccd1 vccd1 _15279_/A sky130_fd_sc_hd__mux2_1
X_17017_ _19413_/Q _16673_/X _17025_/S vssd1 vssd1 vccd1 vccd1 _17018_/A sky130_fd_sc_hd__mux2_1
X_14229_ _13795_/A _14226_/Y _14228_/X vssd1 vssd1 vccd1 vccd1 _14229_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_98_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10338__A2 _19098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17671__A0 _19671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17075__S _17075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _09783_/A vssd1 vssd1 vccd1 vccd1 _09770_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12801__A _13042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18968_ _19589_/CLK _18968_/D vssd1 vssd1 vccd1 vccd1 _18968_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17919_ _19811_/Q _19813_/Q _19812_/Q _18070_/A vssd1 vssd1 vccd1 vccd1 _18079_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_113_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18899_ _19165_/CLK _18899_/D vssd1 vssd1 vccd1 vccd1 _18899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17803__S _17805_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14788__A1 _13086_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13460__A1 _13110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10274__B2 _18442_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12248__A _19681_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ _10022_/A vssd1 vssd1 vccd1 vccd1 _09861_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13212__B2 _18625_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09135_ _09135_/A vssd1 vssd1 vccd1 vccd1 _09854_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_147_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10121__S1 _09147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__A1 _12466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11774__B2 _14575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09557__A _09640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09719__A1 _09689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14712__A1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17774__A _17774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14712__B2 _14711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09968_ _19619_/Q _19457_/Q _18903_/Q _18673_/Q _09872_/S _09936_/X vssd1 vssd1 vccd1
+ vccd1 _09969_/B sky130_fd_sc_hd__mux4_1
XFILLER_131_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13279__B2 _18632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12711__A _18630_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09899_ _11147_/A _11151_/A _11150_/A vssd1 vssd1 vccd1 vccd1 _09899_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10188__S1 _09723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11930_ _12408_/A _11930_/B vssd1 vssd1 vccd1 vccd1 _11930_/Y sky130_fd_sc_hd__nor2_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10231__A _10245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14779__A1 _14777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _19735_/Q _11705_/X _11854_/X _11860_/Y vssd1 vssd1 vccd1 vccd1 _17868_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16329__S _16329_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14638__A _14638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _12011_/A _14192_/B _13681_/S vssd1 vssd1 vccd1 vccd1 _13600_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15233__S _15233_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _18590_/Q _19279_/Q _11028_/S vssd1 vssd1 vccd1 vccd1 _10813_/B sky130_fd_sc_hd__mux2_1
XANTENNA__13542__A _13542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _14580_/A _14580_/B vssd1 vssd1 vccd1 vccd1 _14580_/X sky130_fd_sc_hd__or2_1
XFILLER_32_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13451__A1 _13112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11792_ _19733_/Q _11792_/B vssd1 vssd1 vccd1 vccd1 _12117_/B sky130_fd_sc_hd__and2_1
XFILLER_25_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13531_ _18416_/Q _12692_/X _13542_/A _13530_/X vssd1 vssd1 vccd1 vccd1 _18416_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10743_ _10735_/Y _10741_/X _10742_/X _10752_/A vssd1 vssd1 vccd1 vccd1 _10743_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16250_ _16250_/A vssd1 vssd1 vccd1 vccd1 _19098_/D sky130_fd_sc_hd__clkbuf_1
X_13462_ _18391_/Q _13230_/X _13464_/S vssd1 vssd1 vccd1 vccd1 _13463_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10674_ _18760_/Q _18989_/Q _18920_/Q _19218_/Q _10733_/S _10548_/A vssd1 vssd1 vccd1
+ vccd1 _10675_/B sky130_fd_sc_hd__mux4_1
XFILLER_167_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15201_ _18670_/Q _15200_/X _15201_/S vssd1 vssd1 vccd1 vccd1 _15202_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11997__A _11997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12413_ _11979_/A _12408_/Y _12411_/X _12412_/X _11790_/A vssd1 vssd1 vccd1 vccd1
+ _12413_/X sky130_fd_sc_hd__o311a_1
X_16181_ _16093_/X _19064_/Q _16183_/S vssd1 vssd1 vccd1 vccd1 _16182_/A sky130_fd_sc_hd__mux2_1
X_13393_ _19497_/Q _12741_/X _13391_/X _13392_/X vssd1 vssd1 vccd1 vccd1 _13393_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_127_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_154_clock clkbuf_opt_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19633_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__12962__B1 _17882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15132_ _18650_/Q _13873_/X _15111_/A _11205_/A vssd1 vssd1 vccd1 vccd1 _18650_/D
+ sky130_fd_sc_hd__a22o_1
X_12344_ _12344_/A vssd1 vssd1 vccd1 vccd1 _13525_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16999__S _17003_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15900__A0 _14808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15063_ input24/X _14924_/X _14925_/X vssd1 vssd1 vccd1 vccd1 _15063_/X sky130_fd_sc_hd__a21o_1
X_12275_ _12320_/C _12274_/Y _11928_/X vssd1 vssd1 vccd1 vccd1 _12275_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09805__S1 _09875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14014_ _11846_/Y _13730_/X _14013_/X vssd1 vssd1 vccd1 vccd1 _14014_/X sky130_fd_sc_hd__a21bo_1
X_11226_ _11225_/B _11225_/C _11225_/A vssd1 vssd1 vccd1 vccd1 _11226_/Y sky130_fd_sc_hd__a21oi_1
X_19871_ _19871_/CLK _19871_/D vssd1 vssd1 vccd1 vccd1 _19871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_169_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19635_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__15259__A2 _17149_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17653__A0 _19668_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18822_ _19540_/CLK _18822_/D vssd1 vssd1 vccd1 vccd1 _18822_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15408__S _15410_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11157_ _18877_/Q _19335_/Q _11157_/S vssd1 vssd1 vccd1 vccd1 _11157_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10108_ _18836_/Q _19390_/Q _19552_/Q _18804_/Q _10094_/X _10103_/X vssd1 vssd1 vccd1
+ vccd1 _10108_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09569__S0 _09553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18753_ _19696_/CLK _18753_/D vssd1 vssd1 vccd1 vccd1 _18753_/Q sky130_fd_sc_hd__dfxtp_1
X_11088_ _18862_/Q _19320_/Q _11088_/S vssd1 vssd1 vccd1 vccd1 _11088_/X sky130_fd_sc_hd__mux2_1
X_15965_ _15965_/A vssd1 vssd1 vccd1 vccd1 _18982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17405__A0 _16761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17704_ _12617_/B _17703_/Y _17734_/S vssd1 vssd1 vccd1 vccd1 _17704_/X sky130_fd_sc_hd__mux2_1
X_10039_ _09385_/A _10038_/X _09319_/A vssd1 vssd1 vccd1 vccd1 _10039_/X sky130_fd_sc_hd__o21a_1
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14916_ _14711_/X _14914_/X _14915_/Y vssd1 vssd1 vccd1 vccd1 _16696_/A sky130_fd_sc_hd__a21oi_4
X_18684_ _19472_/CLK _18684_/D vssd1 vssd1 vccd1 vccd1 _18684_/Q sky130_fd_sc_hd__dfxtp_1
X_15896_ _14782_/X _18951_/Q _15902_/S vssd1 vssd1 vccd1 vccd1 _15897_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17635_ _17693_/A vssd1 vssd1 vccd1 vccd1 _17658_/S sky130_fd_sc_hd__clkbuf_2
X_14847_ _16781_/A vssd1 vssd1 vccd1 vccd1 _14847_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17566_ _19642_/Q _16787_/A _17568_/S vssd1 vssd1 vccd1 vccd1 _17567_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_107_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19755_/CLK sky130_fd_sc_hd__clkbuf_16
X_14778_ _14825_/A vssd1 vssd1 vccd1 vccd1 _14893_/A sky130_fd_sc_hd__buf_2
X_19305_ _19642_/CLK _19305_/D vssd1 vssd1 vccd1 vccd1 _19305_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13171__B _18623_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16517_ _19216_/Q _15506_/X _16525_/S vssd1 vssd1 vccd1 vccd1 _16518_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13729_ _13922_/A _13729_/B vssd1 vssd1 vccd1 vccd1 _14102_/A sky130_fd_sc_hd__and2b_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17497_ _17497_/A vssd1 vssd1 vccd1 vccd1 _19611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19236_ _19556_/CLK _19236_/D vssd1 vssd1 vccd1 vccd1 _19236_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15195__A1 _15194_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16448_ _16448_/A vssd1 vssd1 vccd1 vccd1 _19185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09949__A1 _09415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19167_ _19553_/CLK _19167_/D vssd1 vssd1 vccd1 vccd1 _19167_/Q sky130_fd_sc_hd__dfxtp_1
X_16379_ _16379_/A vssd1 vssd1 vccd1 vccd1 _19155_/D sky130_fd_sc_hd__clkbuf_1
X_18118_ _18119_/B _18119_/C _19827_/Q vssd1 vssd1 vccd1 vccd1 _18120_/B sky130_fd_sc_hd__a21oi_1
X_19098_ _19612_/CLK _19098_/D vssd1 vssd1 vccd1 vccd1 _19098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18049_ _18051_/B _18051_/C _18039_/X vssd1 vssd1 vccd1 vccd1 _18049_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_174_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15318__S _15322_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09822_ _10055_/S vssd1 vssd1 vccd1 vccd1 _09865_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09753_ _11222_/A _12500_/A vssd1 vssd1 vccd1 vccd1 _09756_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17533__S _17533_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12054__A1_N _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09684_ _09621_/A _09671_/Y _09677_/X _09683_/Y _09394_/A vssd1 vssd1 vccd1 vccd1
+ _09684_/X sky130_fd_sc_hd__o311a_1
XANTENNA__10051__A _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09840__A _11148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09980__S0 _09782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16673__A _16673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_71_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19618_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09118_ _11471_/A _11585_/A _11376_/C _11495_/B vssd1 vssd1 vccd1 vccd1 _09119_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_135_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10390_ _10390_/A _10390_/B vssd1 vssd1 vccd1 vccd1 _10390_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12425__B _14324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_86_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19788_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12060_ _12060_/A vssd1 vssd1 vccd1 vccd1 _12177_/A sky130_fd_sc_hd__buf_2
XANTENNA__15736__B _17463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11011_ _11062_/A _11008_/X _11010_/X _10728_/A vssd1 vssd1 vccd1 vccd1 _11012_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09573__C1 _09247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15110__A1 _18633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15110__B2 _10412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16848__A _16904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12160__B _13598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12962_ _18298_/Q _18297_/Q _12959_/B _17882_/A vssd1 vssd1 vccd1 vccd1 _12962_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _14772_/X _18886_/Q _15758_/S vssd1 vssd1 vccd1 vccd1 _15751_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input10_A io_dbus_rdata[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ _11913_/A _14045_/A vssd1 vssd1 vccd1 vccd1 _11913_/Y sky130_fd_sc_hd__nor2_1
X_14701_ _14802_/B vssd1 vssd1 vccd1 vccd1 _14701_/Y sky130_fd_sc_hd__inv_2
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19613_/CLK sky130_fd_sc_hd__clkbuf_16
X_12893_ _18277_/Q _12895_/C _12893_/C vssd1 vssd1 vccd1 vccd1 _12894_/C sky130_fd_sc_hd__and3_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15681_ _15681_/A vssd1 vssd1 vccd1 vccd1 _18855_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16059__S _16065_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _16784_/X _19577_/Q _17424_/S vssd1 vssd1 vccd1 vccd1 _17421_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _14632_/A vssd1 vssd1 vccd1 vccd1 _18564_/D sky130_fd_sc_hd__clkbuf_1
X_11844_ _11813_/B _11844_/B vssd1 vssd1 vccd1 vccd1 _11844_/X sky130_fd_sc_hd__and2b_1
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15898__S _15902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _18574_/Q _14526_/B _14562_/Y _14560_/X vssd1 vssd1 vccd1 vccd1 _18542_/D
+ sky130_fd_sc_hd__o211a_1
X_17351_ _17351_/A vssd1 vssd1 vccd1 vccd1 _19546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _11836_/B vssd1 vssd1 vccd1 vccd1 _13939_/B sky130_fd_sc_hd__buf_2
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16302_/A vssd1 vssd1 vccd1 vccd1 _19121_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ _14516_/S vssd1 vssd1 vccd1 vccd1 _14589_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_39_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19724_/CLK sky130_fd_sc_hd__clkbuf_16
X_10726_ _10772_/A vssd1 vssd1 vccd1 vccd1 _10726_/X sky130_fd_sc_hd__clkbuf_4
X_14494_ _18517_/Q _12361_/A _14498_/S vssd1 vssd1 vccd1 vccd1 _14495_/A sky130_fd_sc_hd__mux2_1
X_17282_ _17304_/A vssd1 vssd1 vccd1 vccd1 _17291_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_13_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_clock clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_13_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19021_ _19634_/CLK _19021_/D vssd1 vssd1 vccd1 vccd1 _19021_/Q sky130_fd_sc_hd__dfxtp_1
X_13445_ _18383_/Q _13136_/X _13453_/S vssd1 vssd1 vccd1 vccd1 _13446_/A sky130_fd_sc_hd__mux2_1
X_16233_ _16061_/X _19091_/Q _16235_/S vssd1 vssd1 vccd1 vccd1 _16234_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10657_ _09517_/A _10645_/Y _10652_/X _10656_/Y _09392_/A vssd1 vssd1 vccd1 vccd1
+ _10657_/X sky130_fd_sc_hd__o311a_1
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13376_ _13297_/X _13368_/Y _13375_/X _13306_/X _18645_/Q vssd1 vssd1 vccd1 vccd1
+ _13376_/X sky130_fd_sc_hd__a32o_2
X_16164_ _16067_/X _19056_/Q _16172_/S vssd1 vssd1 vccd1 vccd1 _16165_/A sky130_fd_sc_hd__mux2_1
X_10588_ _10593_/A _10585_/X _10587_/X _09517_/A vssd1 vssd1 vccd1 vccd1 _10589_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_86_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12335__B _19754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12327_ _14274_/B _12327_/B vssd1 vssd1 vccd1 vccd1 _12330_/A sky130_fd_sc_hd__xor2_4
X_15115_ _18637_/Q _15109_/X _15111_/X _10196_/A vssd1 vssd1 vccd1 vccd1 _18637_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10410__B2 _10409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16095_ _16095_/A vssd1 vssd1 vccd1 vccd1 _19032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15046_ _15046_/A vssd1 vssd1 vccd1 vccd1 _18614_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12258_ _14241_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _12262_/A sky130_fd_sc_hd__xnor2_4
XFILLER_170_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09564__C1 _09133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ _11317_/A _11325_/C vssd1 vssd1 vccd1 vccd1 _13526_/B sky130_fd_sc_hd__nand2_2
X_19854_ _19855_/CLK _19854_/D vssd1 vssd1 vccd1 vccd1 _19854_/Q sky130_fd_sc_hd__dfxtp_1
X_12189_ _12408_/A vssd1 vssd1 vccd1 vccd1 _12452_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_110_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11910__A1 _19737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18805_ _19326_/CLK _18805_/D vssd1 vssd1 vccd1 vccd1 _18805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15101__A1 _18627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19785_ _19795_/CLK _19785_/D vssd1 vssd1 vccd1 vccd1 _19785_/Q sky130_fd_sc_hd__dfxtp_1
X_16997_ _19404_/Q _16645_/X _17003_/S vssd1 vssd1 vccd1 vccd1 _16998_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18736_ _19714_/CLK _18736_/D vssd1 vssd1 vccd1 vccd1 _18736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15948_ _15066_/X _18975_/Q _15950_/S vssd1 vssd1 vccd1 vccd1 _15949_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14860__B1 _14859_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10021__S0 _10075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18667_ _19452_/CLK _18667_/D vssd1 vssd1 vccd1 vccd1 _18667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15879_ _15879_/A vssd1 vssd1 vccd1 vccd1 _18944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17618_ _15258_/X _17617_/Y _17149_/Y vssd1 vssd1 vccd1 vccd1 _17618_/X sky130_fd_sc_hd__a21o_1
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18598_ _19513_/CLK _18598_/D vssd1 vssd1 vccd1 vccd1 _18598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10410__A1_N _18440_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17549_ _19634_/Q _16761_/A _17557_/S vssd1 vssd1 vccd1 vccd1 _17550_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15601__S _15603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19219_ _19541_/CLK _19219_/D vssd1 vssd1 vccd1 vccd1 _19219_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14915__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12526__A _12526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10937__C1 _09407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14143__A2 _14138_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12154__B2 _12488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12261__A _12286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09805_ _19525_/Q _19139_/Q _19589_/Q _18745_/Q _09803_/X _09875_/A vssd1 vssd1 vccd1
+ vccd1 _09806_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13076__B _18626_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_A io_dbus_rdata[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17263__S _17269_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09736_ _09736_/A vssd1 vssd1 vccd1 vccd1 _10186_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10468__A1 _09554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09667_ _19656_/Q _19073_/Q _19110_/Q _18716_/Q _09600_/A _10280_/A vssd1 vssd1 vccd1
+ vccd1 _09667_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14188__A _14192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13406__A1 _19688_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ _10389_/S vssd1 vssd1 vccd1 vccd1 _10279_/S sky130_fd_sc_hd__clkbuf_4
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09705__S0 _09545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11560_ _12072_/A vssd1 vssd1 vccd1 vccd1 _11560_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10511_ _18596_/Q _19285_/Q _10511_/S vssd1 vssd1 vccd1 vccd1 _10511_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11491_ _18584_/Q vssd1 vssd1 vccd1 vccd1 _14587_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_137_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13230_ _13217_/X _13218_/Y _13228_/X _13229_/X _18627_/Q vssd1 vssd1 vccd1 vccd1
+ _13230_/X sky130_fd_sc_hd__a32o_4
XFILLER_108_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10442_ _10442_/A _10442_/B vssd1 vssd1 vccd1 vccd1 _10442_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13161_ _19858_/Q _12651_/X _12528_/X _18119_/B _13160_/X vssd1 vssd1 vccd1 vccd1
+ _13161_/X sky130_fd_sc_hd__a221o_1
XFILLER_137_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17438__S _17446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10373_ _10373_/A _10373_/B _10373_/C vssd1 vssd1 vccd1 vccd1 _10373_/X sky130_fd_sc_hd__or3_4
XFILLER_152_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14651__A _14654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12112_ _12112_/A _12112_/B vssd1 vssd1 vccd1 vccd1 _12114_/A sky130_fd_sc_hd__nor2_2
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input58_A io_ibus_inst[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ _13110_/A _18342_/Q _13092_/S vssd1 vssd1 vccd1 vccd1 _13093_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12043_ _12043_/A _12067_/D vssd1 vssd1 vccd1 vccd1 _12044_/B sky130_fd_sc_hd__nand2_1
X_16920_ _17319_/B _16920_/B vssd1 vssd1 vccd1 vccd1 _16977_/A sky130_fd_sc_hd__nand2_4
XFILLER_172_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16851_ _16851_/A vssd1 vssd1 vccd1 vccd1 _19339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15802_ _15055_/X _18910_/Q _15802_/S vssd1 vssd1 vccd1 vccd1 _15803_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19570_ _19636_/CLK _19570_/D vssd1 vssd1 vccd1 vccd1 _19570_/Q sky130_fd_sc_hd__dfxtp_1
X_16782_ _16781_/X _19318_/Q _16791_/S vssd1 vssd1 vccd1 vccd1 _16783_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13994_ _13997_/S _13885_/X _13993_/X vssd1 vssd1 vccd1 vccd1 _13994_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09480__A _09480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18521_ _19079_/CLK _18521_/D vssd1 vssd1 vccd1 vccd1 _18521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ _15733_/A vssd1 vssd1 vccd1 vccd1 _18879_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10459__B2 _10458_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ _18292_/Q _12945_/B vssd1 vssd1 vccd1 vccd1 _12947_/B sky130_fd_sc_hd__nor2_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09864__A3 _09863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11515__A _18575_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18452_ _19692_/CLK _18452_/D vssd1 vssd1 vccd1 vccd1 _18452_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_122_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _16744_/A _17535_/B vssd1 vssd1 vccd1 vccd1 _15721_/A sky130_fd_sc_hd__nor2_2
X_12876_ _12885_/D vssd1 vssd1 vccd1 vccd1 _12883_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _17403_/A vssd1 vssd1 vccd1 vccd1 _19569_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14615_ _14624_/A _14615_/B vssd1 vssd1 vccd1 vccd1 _14616_/A sky130_fd_sc_hd__and2_1
XFILLER_159_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18383_ _19780_/CLK _18383_/D vssd1 vssd1 vccd1 vccd1 _18383_/Q sky130_fd_sc_hd__dfxtp_1
X_11827_ _18356_/Q _11827_/B vssd1 vssd1 vccd1 vccd1 _11827_/X sky130_fd_sc_hd__and2_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15595_ _18817_/Q _15487_/X _15603_/S vssd1 vssd1 vccd1 vccd1 _15596_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17334_/A vssd1 vssd1 vccd1 vccd1 _19538_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _11888_/C vssd1 vssd1 vccd1 vccd1 _11758_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14546_ _18535_/Q _14522_/X _14545_/Y _14535_/X vssd1 vssd1 vccd1 vccd1 _18535_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ _10805_/A vssd1 vssd1 vccd1 vccd1 _10710_/A sky130_fd_sc_hd__clkbuf_4
X_17265_ _19508_/Q _16664_/X _17269_/S vssd1 vssd1 vccd1 vccd1 _17266_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11689_ _11776_/A _13996_/A vssd1 vssd1 vccd1 vccd1 _11695_/A sky130_fd_sc_hd__or2_1
X_14477_ _14477_/A vssd1 vssd1 vccd1 vccd1 _18509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19004_ _19555_/CLK _19004_/D vssd1 vssd1 vccd1 vccd1 _19004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16216_ _16033_/X _19083_/Q _16224_/S vssd1 vssd1 vccd1 vccd1 _16217_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13428_ _18414_/Q _13428_/B vssd1 vssd1 vccd1 vccd1 _13428_/X sky130_fd_sc_hd__and2_1
XFILLER_139_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17196_ _19485_/Q _17195_/X _17206_/S vssd1 vssd1 vccd1 vccd1 _17197_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17348__S _17352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13359_ _19817_/Q vssd1 vssd1 vccd1 vccd1 _18094_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16147_ _16147_/A vssd1 vssd1 vccd1 vccd1 _19048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18033__A _18033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10490__S0 _10450_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16078_ _16077_/X _19027_/Q _16081_/S vssd1 vssd1 vccd1 vccd1 _16079_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_47_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15029_ _18453_/Q _13386_/B _15051_/S vssd1 vssd1 vccd1 vccd1 _15029_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19837_ _19838_/CLK _19837_/D vssd1 vssd1 vccd1 vccd1 _19837_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_111_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15086__A0 _14555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16488__A _16488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16919__C _16919_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19768_ _19859_/CLK _19768_/D vssd1 vssd1 vccd1 vccd1 _19768_/Q sky130_fd_sc_hd__dfxtp_1
Xinput2 io_dbus_rdata[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_2
XANTENNA__13636__A1 _12282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09521_ _10392_/A _09521_/B vssd1 vssd1 vccd1 vccd1 _09521_/Y sky130_fd_sc_hd__nor2_1
X_18719_ _19595_/CLK _18719_/D vssd1 vssd1 vccd1 vccd1 _18719_/Q sky130_fd_sc_hd__dfxtp_1
X_19699_ _19699_/CLK _19699_/D vssd1 vssd1 vccd1 vccd1 _19699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09452_ _09171_/A _09450_/X _09454_/A vssd1 vssd1 vccd1 vccd1 _09452_/X sky130_fd_sc_hd__a21o_1
XFILLER_80_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09383_ _10144_/A vssd1 vssd1 vccd1 vccd1 _10068_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15331__S _15333_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10083__C1 _09230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17258__S _17258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15567__A _16822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12127__B2 _12487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17782__A _17782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09719_ _09689_/X _09712_/X _09714_/X _09718_/X _09248_/A vssd1 vssd1 vccd1 vccd1
+ _09719_/X sky130_fd_sc_hd__a311o_2
X_10991_ _19502_/Q _19116_/Q _19566_/Q _18722_/Q _10668_/A _10960_/X vssd1 vssd1 vccd1
+ vccd1 _10992_/B sky130_fd_sc_hd__mux4_2
XFILLER_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12730_ _18205_/A vssd1 vssd1 vccd1 vccd1 _12731_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _18335_/Q _12810_/A vssd1 vssd1 vccd1 vccd1 _12661_/X sky130_fd_sc_hd__or2_1
XANTENNA__14588__C1 _14585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10861__A1 _10548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _18575_/Q _14553_/A _15095_/B vssd1 vssd1 vccd1 vccd1 _11613_/C sky130_fd_sc_hd__mux2_1
X_14400_ _14400_/A vssd1 vssd1 vccd1 vccd1 _18478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12592_ _12808_/B _12582_/X _12584_/X _19841_/Q _12591_/X vssd1 vssd1 vccd1 vccd1
+ _12592_/X sky130_fd_sc_hd__a221o_2
X_15380_ _18738_/Q _15194_/X _15384_/S vssd1 vssd1 vccd1 vccd1 _15381_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14331_ _14331_/A vssd1 vssd1 vccd1 vccd1 _14331_/Y sky130_fd_sc_hd__inv_2
X_11543_ _15093_/S vssd1 vssd1 vccd1 vccd1 _14032_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12166__A _19678_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11070__A _11070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17050_ _19428_/Q _16721_/X _17058_/S vssd1 vssd1 vccd1 vccd1 _17051_/A sky130_fd_sc_hd__mux2_1
X_14262_ _14262_/A _14265_/B vssd1 vssd1 vccd1 vccd1 _14262_/X sky130_fd_sc_hd__or2_1
XFILLER_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11474_ _11474_/A _11474_/B vssd1 vssd1 vccd1 vccd1 _13584_/A sky130_fd_sc_hd__nor2_1
XFILLER_13_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13213_ _18356_/Q _13246_/B vssd1 vssd1 vccd1 vccd1 _13213_/X sky130_fd_sc_hd__or2_1
XFILLER_7_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16001_ _14918_/X _18999_/Q _16005_/S vssd1 vssd1 vccd1 vccd1 _16002_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10425_ _10432_/A _10421_/X _10424_/X _09459_/X vssd1 vssd1 vccd1 vccd1 _10425_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16072__S _16081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14193_ _14078_/A _14188_/Y _14192_/Y vssd1 vssd1 vccd1 vccd1 _14193_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_152_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10377__B1 _09434_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13144_ _19793_/Q vssd1 vssd1 vccd1 vccd1 _18023_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10356_ _19257_/Q _19028_/Q _18959_/Q _19353_/Q _11087_/S _09142_/A vssd1 vssd1 vccd1
+ vccd1 _10356_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output164_A _17907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14512__C1 _13401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17952_ _17954_/B _17954_/C _17951_/Y vssd1 vssd1 vccd1 vccd1 _19768_/D sky130_fd_sc_hd__o21a_1
X_13075_ _18110_/B _18110_/C _13074_/Y vssd1 vssd1 vccd1 vccd1 _18334_/D sky130_fd_sc_hd__o21a_1
XFILLER_140_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10287_ _19517_/Q _19131_/Q _19581_/Q _18737_/Q _09342_/A _11113_/A vssd1 vssd1 vccd1
+ vccd1 _10288_/B sky130_fd_sc_hd__mux4_1
X_16903_ _16903_/A vssd1 vssd1 vccd1 vccd1 _19363_/D sky130_fd_sc_hd__clkbuf_1
X_12026_ _12026_/A vssd1 vssd1 vccd1 vccd1 _12026_/X sky130_fd_sc_hd__clkbuf_1
X_17883_ _17883_/A vssd1 vssd1 vccd1 vccd1 _19742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19622_ _19622_/CLK _19622_/D vssd1 vssd1 vccd1 vccd1 _19622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16834_ _16834_/A vssd1 vssd1 vccd1 vccd1 _19334_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13618__A1 _12262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19553_ _19553_/CLK _19553_/D vssd1 vssd1 vccd1 vccd1 _19553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16765_ _16765_/A vssd1 vssd1 vccd1 vccd1 _16765_/X sky130_fd_sc_hd__clkbuf_2
X_13977_ _13977_/A vssd1 vssd1 vccd1 vccd1 _14262_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18504_ _18506_/CLK _18504_/D vssd1 vssd1 vccd1 vccd1 _18504_/Q sky130_fd_sc_hd__dfxtp_2
X_15716_ _15716_/A vssd1 vssd1 vccd1 vccd1 _18871_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12928_ _12897_/B _12933_/D _12927_/Y _12802_/X vssd1 vssd1 vccd1 vccd1 _18286_/D
+ sky130_fd_sc_hd__a211oi_1
X_19484_ _19682_/CLK _19484_/D vssd1 vssd1 vccd1 vccd1 _19484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16696_ _16696_/A vssd1 vssd1 vccd1 vccd1 _16696_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18435_ _18818_/CLK _18435_/D vssd1 vssd1 vccd1 vccd1 _18435_/Q sky130_fd_sc_hd__dfxtp_4
X_15647_ _18841_/Q _15567_/X _15647_/S vssd1 vssd1 vccd1 vccd1 _15648_/A sky130_fd_sc_hd__mux2_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12859_ _12863_/B _12863_/C _12817_/X vssd1 vssd1 vccd1 vccd1 _12859_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18366_ _18402_/CLK _18366_/D vssd1 vssd1 vccd1 vccd1 _18366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15578_ _18812_/Q _15577_/X _15584_/S vssd1 vssd1 vccd1 vccd1 _15579_/A sky130_fd_sc_hd__mux2_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17317_ _19532_/Q _16740_/X _17317_/S vssd1 vssd1 vccd1 vccd1 _17318_/A sky130_fd_sc_hd__mux2_1
X_14529_ _16138_/A _14582_/B vssd1 vssd1 vccd1 vccd1 _14529_/Y sky130_fd_sc_hd__nand2_1
X_18297_ _18402_/CLK _18297_/D vssd1 vssd1 vccd1 vccd1 _18297_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09470__A1 _09434_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17248_ _17304_/A vssd1 vssd1 vccd1 vccd1 _17317_/S sky130_fd_sc_hd__buf_8
XFILLER_128_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17179_ _19480_/Q _17178_/X _17189_/S vssd1 vssd1 vccd1 vccd1 _17180_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10463__S0 _09631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10383__A3 _10382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16710__S _16719_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11139__B _12488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13609__A1 _14168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14282__A1 _14281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11155__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09504_ _10227_/A vssd1 vssd1 vccd1 vccd1 _10400_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09435_ _19691_/Q vssd1 vssd1 vccd1 vccd1 _10905_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_52_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12045__A0 _12041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09366_ _09421_/A _09366_/B vssd1 vssd1 vccd1 vccd1 _09366_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09461__A1 _09434_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ _14570_/A _14716_/A _16138_/B _11516_/A vssd1 vssd1 vccd1 vccd1 _09303_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_119_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12714__A _13108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10210_ _10210_/A _10210_/B vssd1 vssd1 vccd1 vccd1 _10210_/X sky130_fd_sc_hd__or2_1
XFILLER_134_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11020__A1 _10807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ _09723_/X _11187_/Y _11189_/Y _10325_/A vssd1 vssd1 vccd1 vccd1 _11190_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10454__S0 _10401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13529__B _13529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10141_ _19648_/Q _19065_/Q _19102_/Q _18708_/Q _09734_/X _10186_/A vssd1 vssd1 vccd1
+ vccd1 _10141_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17039__A1 _16705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_0_0_clock clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_0_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10072_ _09927_/X _10062_/X _10071_/X _09309_/A _18446_/Q vssd1 vssd1 vccd1 vccd1
+ _12489_/C sky130_fd_sc_hd__a32o_4
XFILLER_0_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13900_ _13918_/S _13898_/X _13899_/X vssd1 vssd1 vccd1 vccd1 _13901_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__15236__S _15239_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14880_ _14879_/X _18600_/Q _14880_/S vssd1 vssd1 vccd1 vccd1 _14881_/A sky130_fd_sc_hd__mux2_1
X_13831_ _13950_/A vssd1 vssd1 vccd1 vccd1 _13832_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14273__A1 _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17451__S _17457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15760__A _15806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16550_ _19231_/Q _15554_/X _16558_/S vssd1 vssd1 vccd1 vccd1 _16551_/A sky130_fd_sc_hd__mux2_1
X_10974_ _18756_/Q _18985_/Q _18916_/Q _19214_/Q _10668_/A _10906_/A vssd1 vssd1 vccd1
+ vccd1 _10975_/B sky130_fd_sc_hd__mux4_1
X_13762_ _13999_/S vssd1 vssd1 vccd1 vccd1 _13918_/S sky130_fd_sc_hd__clkbuf_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15501_ _18788_/Q _15500_/X _15504_/S vssd1 vssd1 vccd1 vccd1 _15502_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10295__C1 _09402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12713_ _12600_/X _12701_/Y _12711_/X _12712_/X _18630_/Q vssd1 vssd1 vccd1 vccd1
+ _12713_/X sky130_fd_sc_hd__a32o_4
X_16481_ _16481_/A vssd1 vssd1 vccd1 vccd1 _19200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13693_ _13677_/X _13692_/X _14103_/A vssd1 vssd1 vccd1 vccd1 _13693_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18220_ _19861_/Q _18222_/C _12948_/X vssd1 vssd1 vccd1 vccd1 _18221_/B sky130_fd_sc_hd__o21ai_1
XFILLER_102_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15432_ _15432_/A vssd1 vssd1 vccd1 vccd1 _18759_/D sky130_fd_sc_hd__clkbuf_1
X_12644_ _12669_/A vssd1 vssd1 vccd1 vccd1 _13418_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_31_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18151_ _18159_/A _18156_/C vssd1 vssd1 vccd1 vccd1 _18151_/Y sky130_fd_sc_hd__nor2_1
XFILLER_157_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12575_ _13440_/S vssd1 vssd1 vccd1 vccd1 _12575_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15363_ _15363_/A vssd1 vssd1 vccd1 vccd1 _18730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09452__A1 _09171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17102_ _16797_/X _19451_/Q _17108_/S vssd1 vssd1 vccd1 vccd1 _17103_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14314_ _14314_/A _14314_/B vssd1 vssd1 vccd1 vccd1 _14314_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18082_ _18170_/A vssd1 vssd1 vccd1 vccd1 _18082_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10693__S0 _10770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11526_ _13579_/B _11526_/B _13587_/A vssd1 vssd1 vccd1 vccd1 _11539_/B sky130_fd_sc_hd__and3b_1
X_15294_ _18700_/Q _15175_/X _15300_/S vssd1 vssd1 vccd1 vccd1 _15295_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17033_ _17033_/A vssd1 vssd1 vccd1 vccd1 _19420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14245_ _13823_/A _14020_/X _14244_/X _14115_/X vssd1 vssd1 vccd1 vccd1 _14245_/X
+ sky130_fd_sc_hd__a211o_1
X_11457_ _11457_/A vssd1 vssd1 vccd1 vccd1 _19079_/D sky130_fd_sc_hd__clkbuf_1
X_10408_ _09411_/A _10400_/Y _10403_/Y _10405_/Y _10407_/Y vssd1 vssd1 vccd1 vccd1
+ _10408_/X sky130_fd_sc_hd__o32a_1
X_14176_ _14178_/B _14176_/B vssd1 vssd1 vccd1 vccd1 _14180_/B sky130_fd_sc_hd__and2_1
X_11388_ _18423_/Q _14802_/B _18421_/Q vssd1 vssd1 vccd1 vccd1 _11388_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_output89_A _12290_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13127_ _13127_/A vssd1 vssd1 vccd1 vccd1 _13127_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10339_ _10327_/A _10338_/X _09616_/A vssd1 vssd1 vccd1 vccd1 _10339_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_140_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18984_ _19698_/CLK _18984_/D vssd1 vssd1 vccd1 vccd1 _18984_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ _17935_/A _17935_/B _17935_/C vssd1 vssd1 vccd1 vccd1 _19763_/D sky130_fd_sc_hd__nor3_1
X_13058_ _18328_/Q _18330_/Q _18329_/Q _13058_/D vssd1 vssd1 vccd1 vccd1 _13069_/D
+ sky130_fd_sc_hd__and4_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12009_ _11130_/A _18503_/Q _12060_/A vssd1 vssd1 vccd1 vccd1 _13595_/A sky130_fd_sc_hd__mux2_4
XFILLER_66_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17866_ _17874_/A _17866_/B vssd1 vssd1 vccd1 vccd1 _17867_/A sky130_fd_sc_hd__or2_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16817_ _16816_/X _19329_/Q _16823_/S vssd1 vssd1 vccd1 vccd1 _16818_/A sky130_fd_sc_hd__mux2_1
X_19605_ _19702_/CLK _19605_/D vssd1 vssd1 vccd1 vccd1 _19605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17797_ _15155_/X _19701_/Q _17805_/S vssd1 vssd1 vccd1 vccd1 _17798_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17361__S _17363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19536_ _19691_/CLK _19536_/D vssd1 vssd1 vccd1 vccd1 _19536_/Q sky130_fd_sc_hd__dfxtp_1
X_16748_ _16748_/A vssd1 vssd1 vccd1 vccd1 _19307_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11406__C _12526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10286__C1 _09393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19467_ _19467_/CLK hold1/X vssd1 vssd1 vccd1 vccd1 _19467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16679_ _16679_/A vssd1 vssd1 vccd1 vccd1 _19286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09220_ _18784_/Q _19013_/Q _18944_/Q _19242_/Q _09190_/A _09149_/A vssd1 vssd1 vccd1
+ vccd1 _09221_/B sky130_fd_sc_hd__mux4_1
XFILLER_146_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18418_ _18578_/CLK _18418_/D vssd1 vssd1 vccd1 vccd1 _18418_/Q sky130_fd_sc_hd__dfxtp_1
X_19398_ _19643_/CLK _19398_/D vssd1 vssd1 vccd1 vccd1 _19398_/Q sky130_fd_sc_hd__dfxtp_1
X_09151_ _11028_/S vssd1 vssd1 vccd1 vccd1 _09152_/A sky130_fd_sc_hd__clkbuf_4
X_18349_ _18386_/CLK _18349_/D vssd1 vssd1 vccd1 vccd1 _18349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09082_ _09088_/A vssd1 vssd1 vccd1 vccd1 _11358_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput60 io_ibus_inst[4] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_1
Xinput71 io_irq_uart_irq vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10987__S1 _10739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16440__S _16442_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09984_ _09984_/A vssd1 vssd1 vccd1 vccd1 _09984_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_89_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15056__S _15056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12266__B1 _19751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11069__B2 _12458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09682__A1 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_169_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10911__S1 _10910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09418_ _18848_/Q _19402_/Q _19564_/Q _18816_/Q _09367_/S _09364_/A vssd1 vssd1 vccd1
+ vccd1 _09419_/B sky130_fd_sc_hd__mux4_1
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10690_ _10683_/X _10685_/X _10687_/X _10689_/X _09244_/A vssd1 vssd1 vccd1 vccd1
+ _10690_/X sky130_fd_sc_hd__a221o_2
X_09349_ _09367_/S vssd1 vssd1 vccd1 vccd1 _09369_/S sky130_fd_sc_hd__buf_2
XFILLER_8_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10229__A _11119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12360_ _12361_/A _12387_/C vssd1 vssd1 vccd1 vccd1 _12362_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11311_ _11528_/A _11310_/X _11564_/A vssd1 vssd1 vccd1 vccd1 _11592_/A sky130_fd_sc_hd__o21bai_2
XFILLER_166_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12291_ _19752_/Q _12292_/B vssd1 vssd1 vccd1 vccd1 _12293_/A sky130_fd_sc_hd__nor2_1
XFILLER_107_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14030_ _13931_/A _14019_/X _14029_/X _13871_/X vssd1 vssd1 vccd1 vccd1 _14030_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11242_ _11242_/A _11242_/B _11242_/C vssd1 vssd1 vccd1 vccd1 _11242_/Y sky130_fd_sc_hd__nand3_1
XFILLER_107_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17446__S _17446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11173_ _09689_/X _11166_/X _11168_/X _11172_/X _09248_/A vssd1 vssd1 vccd1 vccd1
+ _11173_/X sky130_fd_sc_hd__a311o_4
XFILLER_164_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18131__A _19830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18209__B1 _12948_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input40_A io_ibus_inst[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ _09278_/A _10112_/X _10123_/X _09285_/A _18445_/Q vssd1 vssd1 vccd1 vccd1
+ _11139_/A sky130_fd_sc_hd__a32o_4
XANTENNA__09753__A _11222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15981_ _14808_/X _18990_/Q _15983_/S vssd1 vssd1 vccd1 vccd1 _15982_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14494__A1 _12361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17720_ _18478_/Q _18479_/Q _17720_/C vssd1 vssd1 vccd1 vccd1 _17728_/B sky130_fd_sc_hd__or3_1
X_10055_ _18606_/Q _19295_/Q _10055_/S vssd1 vssd1 vccd1 vccd1 _10055_/X sky130_fd_sc_hd__mux2_1
X_14932_ _18476_/Q _18477_/Q _14932_/C vssd1 vssd1 vccd1 vccd1 _14955_/C sky130_fd_sc_hd__and3_1
XFILLER_169_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17651_ _17656_/B _17651_/B vssd1 vssd1 vccd1 vccd1 _17651_/Y sky130_fd_sc_hd__nand2_2
XFILLER_76_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14863_ _14871_/B _14945_/B _14863_/C vssd1 vssd1 vccd1 vccd1 _14863_/X sky130_fd_sc_hd__and3b_1
XFILLER_169_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14246__A1 _12265_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10411__B _12482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16602_ _16602_/A vssd1 vssd1 vccd1 vccd1 _19256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13814_ _13965_/S _13812_/X _13813_/Y vssd1 vssd1 vccd1 vccd1 _13814_/Y sky130_fd_sc_hd__a21boi_1
X_17582_ _19649_/Q _16809_/A _17590_/S vssd1 vssd1 vccd1 vccd1 _17583_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14794_ _14794_/A vssd1 vssd1 vccd1 vccd1 _18593_/D sky130_fd_sc_hd__clkbuf_1
X_19321_ _19513_/CLK _19321_/D vssd1 vssd1 vccd1 vccd1 _19321_/Q sky130_fd_sc_hd__dfxtp_1
X_16533_ _16533_/A vssd1 vssd1 vccd1 vccd1 _19223_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13745_ _13881_/S vssd1 vssd1 vccd1 vccd1 _13745_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10957_ _19600_/Q _19438_/Q _18884_/Q _18654_/Q _10909_/X _10910_/X vssd1 vssd1 vccd1
+ vccd1 _10958_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10838__S _10886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12009__A0 _11130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19252_ _19726_/CLK _19252_/D vssd1 vssd1 vccd1 vccd1 _19252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16464_ _16080_/X _19193_/Q _16464_/S vssd1 vssd1 vccd1 vccd1 _16465_/A sky130_fd_sc_hd__mux2_1
X_13676_ _13845_/S vssd1 vssd1 vccd1 vccd1 _13965_/S sky130_fd_sc_hd__clkbuf_2
X_10888_ _09353_/A _10885_/Y _10887_/Y _10701_/A vssd1 vssd1 vccd1 vccd1 _10888_/X
+ sky130_fd_sc_hd__o211a_1
X_18203_ _19855_/Q _18201_/B _18170_/X vssd1 vssd1 vccd1 vccd1 _18203_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12338__B _13529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15415_ _16503_/B _17535_/B vssd1 vssd1 vccd1 vccd1 _15472_/A sky130_fd_sc_hd__nor2_2
X_12627_ _18369_/Q _13236_/A _12623_/X _12626_/X vssd1 vssd1 vccd1 vccd1 _12627_/X
+ sky130_fd_sc_hd__a211o_1
X_19183_ _19633_/CLK _19183_/D vssd1 vssd1 vccd1 vccd1 _19183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16395_ _16395_/A vssd1 vssd1 vccd1 vccd1 _19162_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14834__A _15077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18134_ _18142_/D vssd1 vssd1 vccd1 vccd1 _18140_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09928__A _09928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15346_ _15346_/A vssd1 vssd1 vccd1 vccd1 _18722_/D sky130_fd_sc_hd__clkbuf_1
X_12558_ _12712_/A vssd1 vssd1 vccd1 vccd1 _12558_/X sky130_fd_sc_hd__buf_2
XANTENNA__09520__S1 _09483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18065_ _18067_/B _18067_/C _18039_/X vssd1 vssd1 vccd1 vccd1 _18065_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11509_ _18576_/Q vssd1 vssd1 vccd1 vccd1 _14568_/A sky130_fd_sc_hd__buf_2
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15277_ _15277_/A vssd1 vssd1 vccd1 vccd1 _18692_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12489_ _12495_/A _12495_/B _12489_/C vssd1 vssd1 vccd1 vccd1 _12490_/A sky130_fd_sc_hd__and3_1
XANTENNA__09189__B1 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17016_ _17062_/S vssd1 vssd1 vccd1 vccd1 _17025_/S sky130_fd_sc_hd__clkbuf_4
X_14228_ _14142_/A _14223_/Y _14227_/Y _13864_/A vssd1 vssd1 vccd1 vccd1 _14228_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16260__S _16268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14159_ _13832_/A _14145_/B _14012_/X vssd1 vssd1 vccd1 vccd1 _14159_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11091__S0 _10348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09663__A _10245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18967_ _19833_/CLK _18967_/D vssd1 vssd1 vccd1 vccd1 _18967_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14485__A1 _19751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17880__A _17882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17918_ _19809_/Q _19808_/Q _19810_/Q _18062_/A vssd1 vssd1 vccd1 vccd1 _18070_/A
+ sky130_fd_sc_hd__and4_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18898_ _19642_/CLK _18898_/D vssd1 vssd1 vccd1 vccd1 _18898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17849_ _15232_/X _19725_/Q _17849_/S vssd1 vssd1 vccd1 vccd1 _17850_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17091__S _17097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19519_ _19647_/CLK _19519_/D vssd1 vssd1 vccd1 vccd1 _19519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_170_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16934__A0 _16761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09203_ _10074_/A vssd1 vssd1 vccd1 vccd1 _10022_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09134_ _09134_/A vssd1 vssd1 vccd1 vccd1 _09135_/A sky130_fd_sc_hd__buf_2
XANTENNA__09838__A _18450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14712__A2 _14703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16170__S _16172_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_95_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09967_ _09879_/A _09966_/X _09892_/A vssd1 vssd1 vccd1 vccd1 _09967_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12711__B _12711_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14476__A1 _19747_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09898_ _09898_/A _12499_/A vssd1 vssd1 vccd1 vccd1 _11150_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _11857_/Y _11858_/X _11859_/X vssd1 vssd1 vccd1 vccd1 _11860_/Y sky130_fd_sc_hd__o21ai_2
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17178__A0 _18437_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10811_ _09926_/A _10799_/X _10809_/X _09306_/A _10810_/X vssd1 vssd1 vccd1 vccd1
+ _12465_/A sky130_fd_sc_hd__a32oi_4
XFILLER_72_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ _19733_/Q _11792_/B vssd1 vssd1 vccd1 vccd1 _11794_/A sky130_fd_sc_hd__nor2_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11732__A_N _13653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13530_ _13521_/X _13522_/X _13529_/X _14519_/B vssd1 vssd1 vccd1 vccd1 _13530_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10896__S0 _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10742_ _19249_/Q _19020_/Q _18951_/Q _19345_/Q _10669_/A _10670_/X vssd1 vssd1 vccd1
+ vccd1 _10742_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16925__A0 _16749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13461_ _13461_/A vssd1 vssd1 vccd1 vccd1 _18390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10673_ _10665_/Y _10671_/X _10672_/X _10873_/A vssd1 vssd1 vccd1 vccd1 _10673_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16345__S _16351_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14654__A _14654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18126__A _18170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15200_ _16702_/A vssd1 vssd1 vccd1 vccd1 _15200_/X sky130_fd_sc_hd__clkbuf_2
X_12412_ _19688_/Q _12412_/B vssd1 vssd1 vccd1 vccd1 _12412_/X sky130_fd_sc_hd__or2_1
XFILLER_127_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16180_ _16180_/A vssd1 vssd1 vccd1 vccd1 _19063_/D sky130_fd_sc_hd__clkbuf_1
X_13392_ _19687_/Q _13251_/X _12743_/X _18411_/Q vssd1 vssd1 vccd1 vccd1 _13392_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15131_ _18649_/Q _13873_/X _15111_/A _11202_/A vssd1 vssd1 vccd1 vccd1 _18649_/D
+ sky130_fd_sc_hd__a22o_1
X_12343_ _19754_/Q _12186_/X _12339_/X _12342_/Y vssd1 vssd1 vccd1 vccd1 _12343_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_127_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12274_ _18373_/Q _12251_/X _17693_/A vssd1 vssd1 vccd1 vccd1 _12274_/Y sky130_fd_sc_hd__o21ai_1
X_15062_ _14875_/X _15069_/B _15059_/X _15061_/X vssd1 vssd1 vccd1 vccd1 _15062_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_141_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14013_ _13726_/X _13999_/X _14011_/X _14012_/X vssd1 vssd1 vccd1 vccd1 _14013_/X
+ sky130_fd_sc_hd__a211o_1
X_11225_ _11225_/A _11225_/B _11225_/C vssd1 vssd1 vccd1 vccd1 _11225_/X sky130_fd_sc_hd__and3_1
X_19870_ _19871_/CLK _19870_/D vssd1 vssd1 vccd1 vccd1 _19870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11156_ _18614_/Q _19303_/Q _11156_/S vssd1 vssd1 vccd1 vccd1 _11156_/X sky130_fd_sc_hd__mux2_1
X_18821_ _19537_/CLK _18821_/D vssd1 vssd1 vccd1 vccd1 _18821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13717__B _13720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10107_ _10107_/A _10107_/B vssd1 vssd1 vccd1 vccd1 _10107_/X sky130_fd_sc_hd__or2_1
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18752_ _19647_/CLK _18752_/D vssd1 vssd1 vccd1 vccd1 _18752_/Q sky130_fd_sc_hd__dfxtp_1
X_15964_ _14714_/X _18982_/Q _15972_/S vssd1 vssd1 vccd1 vccd1 _15965_/A sky130_fd_sc_hd__mux2_1
X_11087_ _18599_/Q _19288_/Q _11087_/S vssd1 vssd1 vccd1 vccd1 _11087_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09569__S1 _09555_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17703_ _17710_/B _17703_/B vssd1 vssd1 vccd1 vccd1 _17703_/Y sky130_fd_sc_hd__nand2_1
X_10038_ _19424_/Q _19200_/Q _19717_/Q _19168_/Q _09866_/A _09869_/A vssd1 vssd1 vccd1
+ vccd1 _10038_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10489__C1 _09529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14915_ input9/X _14901_/X _14904_/X vssd1 vssd1 vccd1 vccd1 _14915_/Y sky130_fd_sc_hd__a21oi_1
X_18683_ _19472_/CLK _18683_/D vssd1 vssd1 vccd1 vccd1 _18683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09894__A1 _09415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15895_ _15895_/A vssd1 vssd1 vccd1 vccd1 _18950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15424__S _15426_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17634_ _17640_/B _17634_/B vssd1 vssd1 vccd1 vccd1 _17634_/Y sky130_fd_sc_hd__nand2_2
X_14846_ _16677_/A vssd1 vssd1 vccd1 vccd1 _16781_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17565_ _17565_/A vssd1 vssd1 vccd1 vccd1 _19641_/D sky130_fd_sc_hd__clkbuf_1
X_14777_ _18432_/Q _13211_/B _14992_/S vssd1 vssd1 vccd1 vccd1 _14777_/X sky130_fd_sc_hd__mux2_1
X_11989_ _12098_/B vssd1 vssd1 vccd1 vccd1 _11989_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19304_ _19626_/CLK _19304_/D vssd1 vssd1 vccd1 vccd1 _19304_/Q sky130_fd_sc_hd__dfxtp_1
X_16516_ _16573_/S vssd1 vssd1 vccd1 vccd1 _16525_/S sky130_fd_sc_hd__buf_2
XFILLER_44_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13728_ _13594_/X _13696_/X _13870_/B _13727_/X vssd1 vssd1 vccd1 vccd1 _13728_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17496_ _19611_/Q _16686_/X _17496_/S vssd1 vssd1 vccd1 vccd1 _17497_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19235_ _19557_/CLK _19235_/D vssd1 vssd1 vccd1 vccd1 _19235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16447_ _16055_/X _19185_/Q _16453_/S vssd1 vssd1 vccd1 vccd1 _16448_/A sky130_fd_sc_hd__mux2_1
X_13659_ _12282_/A _13658_/X _13659_/S vssd1 vssd1 vccd1 vccd1 _13659_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16255__S _16257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19166_ _19715_/CLK _19166_/D vssd1 vssd1 vccd1 vccd1 _19166_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10639__S0 _10500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16378_ _19155_/Q _15516_/X _16380_/S vssd1 vssd1 vccd1 vccd1 _16379_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18117_ _18119_/B _18119_/C _18116_/Y vssd1 vssd1 vccd1 vccd1 _19826_/D sky130_fd_sc_hd__o21a_1
XFILLER_145_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15329_ _18716_/Q _15226_/X _15333_/S vssd1 vssd1 vccd1 vccd1 _15330_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17341__A0 _16774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19097_ _19579_/CLK _19097_/D vssd1 vssd1 vccd1 vccd1 _19097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18048_ _19801_/Q _18045_/B _18047_/Y vssd1 vssd1 vccd1 vccd1 _19801_/D sky130_fd_sc_hd__o21a_1
XFILLER_145_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_117_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12812__A _18225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09821_ _09821_/A vssd1 vssd1 vccd1 vccd1 _09821_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09393__A _09393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10192__A1 _09621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17814__S _17816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ _09430_/A _09741_/X _09750_/X _09625_/X _09751_/Y vssd1 vssd1 vccd1 vccd1
+ _12500_/A sky130_fd_sc_hd__o32a_4
XFILLER_100_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11837__D_N _13996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09683_ _09671_/A _09678_/X _09682_/X vssd1 vssd1 vccd1 vccd1 _09683_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13643__A _13643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09840__B _12497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19709_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09980__S1 _09979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14630__A1 _18564_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11444__A1 _18343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10652__C1 _10764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13197__B2 _18624_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17785__A _17853_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09117_ _11361_/A vssd1 vssd1 vccd1 vccd1 _11585_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10507__A _11082_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14697__A1 _14589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15894__A0 _14772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14697__B2 input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _18979_/Q _11010_/B vssd1 vssd1 vccd1 vccd1 _11010_/X sky130_fd_sc_hd__or2_1
XFILLER_78_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10802__S0 _10719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12961_ _12961_/A _12961_/B vssd1 vssd1 vccd1 vccd1 _18297_/D sky130_fd_sc_hd__nor2_1
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09876__A1 _09826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _18423_/Q vssd1 vssd1 vccd1 vccd1 _14802_/A sky130_fd_sc_hd__inv_2
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11912_ _12476_/B _11831_/X _11911_/X vssd1 vssd1 vccd1 vccd1 _14059_/B sky130_fd_sc_hd__a21o_2
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11683__A1 _17143_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _18855_/Q _15510_/X _15686_/S vssd1 vssd1 vccd1 vccd1 _15681_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12892_ _12895_/C _12893_/C _18277_/Q vssd1 vssd1 vccd1 vccd1 _12894_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12880__B1 _12869_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _14654_/A _14631_/B vssd1 vssd1 vccd1 vccd1 _14632_/A sky130_fd_sc_hd__and2_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _11843_/A vssd1 vssd1 vccd1 vccd1 _13984_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17350_ _16787_/X _19546_/Q _17352_/S vssd1 vssd1 vccd1 vccd1 _17351_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _14562_/A _14582_/B vssd1 vssd1 vccd1 vccd1 _14562_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11774_ _12466_/A _11831_/A _11911_/C _14575_/A vssd1 vssd1 vccd1 vccd1 _11836_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16301_ _16055_/X _19121_/Q _16307_/S vssd1 vssd1 vccd1 vccd1 _16302_/A sky130_fd_sc_hd__mux2_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _13513_/A vssd1 vssd1 vccd1 vccd1 _18414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10725_ _10725_/A vssd1 vssd1 vccd1 vccd1 _10772_/A sky130_fd_sc_hd__buf_2
X_17281_ _17281_/A vssd1 vssd1 vccd1 vccd1 _19515_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14493_ _14493_/A vssd1 vssd1 vccd1 vccd1 _18516_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16374__A1 _15510_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16075__S _16081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19020_ _19635_/CLK _19020_/D vssd1 vssd1 vccd1 vccd1 _19020_/Q sky130_fd_sc_hd__dfxtp_1
X_16232_ _16232_/A vssd1 vssd1 vccd1 vccd1 _19090_/D sky130_fd_sc_hd__clkbuf_1
X_13444_ _13512_/S vssd1 vssd1 vccd1 vccd1 _13453_/S sky130_fd_sc_hd__buf_2
XFILLER_174_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10656_ _10640_/A _10653_/X _10655_/X vssd1 vssd1 vccd1 vccd1 _10656_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16163_ _16209_/S vssd1 vssd1 vccd1 vccd1 _16172_/S sky130_fd_sc_hd__clkbuf_8
X_13375_ _18645_/Q _15018_/B vssd1 vssd1 vccd1 vccd1 _13375_/X sky130_fd_sc_hd__or2_1
X_10587_ _10640_/A _10587_/B vssd1 vssd1 vccd1 vccd1 _10587_/X sky130_fd_sc_hd__or2_1
XFILLER_6_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15114_ _18636_/Q _15109_/X _15111_/X _11137_/A vssd1 vssd1 vccd1 vccd1 _18636_/D
+ sky130_fd_sc_hd__a22o_1
X_12326_ _12348_/A _14265_/A _12305_/B vssd1 vssd1 vccd1 vccd1 _12327_/B sky130_fd_sc_hd__a21bo_1
XFILLER_127_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16094_ _16093_/X _19032_/Q _16097_/S vssd1 vssd1 vccd1 vccd1 _16095_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09239__S0 _09190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15885__A0 _14729_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15045_ _15044_/X _18614_/Q _15056_/S vssd1 vssd1 vccd1 vccd1 _15046_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12257_ _13567_/A _14227_/A _12230_/B vssd1 vssd1 vccd1 vccd1 _12258_/B sky130_fd_sc_hd__o21a_2
XFILLER_69_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11208_ _11205_/Y _11284_/C _13568_/A vssd1 vssd1 vccd1 vccd1 _11208_/Y sky130_fd_sc_hd__a21oi_1
X_19853_ _19871_/CLK _19853_/D vssd1 vssd1 vccd1 vccd1 _19853_/Q sky130_fd_sc_hd__dfxtp_1
X_12188_ _19748_/Q _12188_/B vssd1 vssd1 vccd1 vccd1 _12188_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_96_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18804_ _19584_/CLK _18804_/D vssd1 vssd1 vccd1 vccd1 _18804_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15101__A2 _13566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ _11139_/A _12488_/A vssd1 vssd1 vccd1 vccd1 _11139_/X sky130_fd_sc_hd__and2_1
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19784_ _19790_/CLK _19784_/D vssd1 vssd1 vccd1 vccd1 _19784_/Q sky130_fd_sc_hd__dfxtp_1
X_16996_ _16996_/A vssd1 vssd1 vccd1 vccd1 _19403_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18735_ _19643_/CLK _18735_/D vssd1 vssd1 vccd1 vccd1 _18735_/Q sky130_fd_sc_hd__dfxtp_1
X_15947_ _15947_/A vssd1 vssd1 vccd1 vccd1 _18974_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14559__A _14559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14860__A1 _18439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10021__S1 _09147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18666_ _19551_/CLK _18666_/D vssd1 vssd1 vccd1 vccd1 _18666_/Q sky130_fd_sc_hd__dfxtp_1
X_15878_ _15076_/X _18944_/Q _15878_/S vssd1 vssd1 vccd1 vccd1 _15879_/A sky130_fd_sc_hd__mux2_1
X_17617_ _17621_/A _17621_/C vssd1 vssd1 vccd1 vccd1 _17617_/Y sky130_fd_sc_hd__xnor2_4
X_14829_ _14840_/B _14829_/B _14829_/C vssd1 vssd1 vccd1 vccd1 _14829_/X sky130_fd_sc_hd__and3b_1
X_18597_ _19414_/CLK _18597_/D vssd1 vssd1 vccd1 vccd1 _18597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17548_ _17605_/S vssd1 vssd1 vccd1 vccd1 _17557_/S sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_43_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10032__A_N _09936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16365__A1 _15497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17479_ _19603_/Q _16661_/X _17485_/S vssd1 vssd1 vccd1 vccd1 _17480_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11711__A _19662_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19218_ _19442_/CLK _19218_/D vssd1 vssd1 vccd1 vccd1 _19218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19149_ _19698_/CLK _19149_/D vssd1 vssd1 vccd1 vccd1 _19149_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16713__S _16719_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15329__S _15333_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13351__A1 _12757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10165__A1 _09996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09650__S0 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09804_ _09810_/A vssd1 vssd1 vccd1 vccd1 _09875_/A sky130_fd_sc_hd__buf_2
XANTENNA__17544__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10260__S1 _09697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09735_ _09735_/A vssd1 vssd1 vccd1 vccd1 _09736_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_153_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19631_/CLK sky130_fd_sc_hd__clkbuf_16
X_09666_ _09732_/A _09666_/B vssd1 vssd1 vccd1 vccd1 _09666_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15999__S _16005_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09597_ _09671_/A vssd1 vssd1 vccd1 vccd1 _10325_/A sky130_fd_sc_hd__buf_2
XFILLER_36_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09705__S1 _10080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_168_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19614_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10510_ _10384_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10510_/X sky130_fd_sc_hd__and2b_1
X_11490_ _18585_/Q vssd1 vssd1 vccd1 vccd1 _14589_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10441_ _19513_/Q _19127_/Q _19577_/Q _18733_/Q _10230_/X _10245_/X vssd1 vssd1 vccd1
+ vccd1 _10442_/B sky130_fd_sc_hd__mux4_1
XFILLER_109_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13590__A1 _12450_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13160_ _13154_/X _13155_/X _13158_/X _12666_/B _17934_/B vssd1 vssd1 vccd1 vccd1
+ _13160_/X sky130_fd_sc_hd__o32a_1
XFILLER_124_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10372_ _10432_/A _10369_/X _10371_/X _09459_/X vssd1 vssd1 vccd1 vccd1 _10373_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12111_ _12111_/A _13608_/A vssd1 vssd1 vccd1 vccd1 _12112_/B sky130_fd_sc_hd__nor2_1
XANTENNA__15239__S _15239_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13091_ _13091_/A vssd1 vssd1 vccd1 vccd1 _18341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12042_ _19742_/Q vssd1 vssd1 vccd1 vccd1 _12067_/B sky130_fd_sc_hd__buf_4
XFILLER_105_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_106_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19759_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_151_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10156__A1 _09984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16850_ _19339_/Q _16639_/X _16858_/S vssd1 vssd1 vccd1 vccd1 _16851_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15801_ _15801_/A vssd1 vssd1 vccd1 vccd1 _18909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09761__A _09978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16781_ _16781_/A vssd1 vssd1 vccd1 vccd1 _16781_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13993_ _13993_/A _13993_/B vssd1 vssd1 vccd1 vccd1 _13993_/X sky130_fd_sc_hd__or2_1
XFILLER_46_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18520_ _19079_/CLK _18520_/D vssd1 vssd1 vccd1 vccd1 _18520_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15732_ _18879_/Q _15586_/X _15734_/S vssd1 vssd1 vccd1 vccd1 _15733_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12944_ _12991_/A vssd1 vssd1 vccd1 vccd1 _12983_/A sky130_fd_sc_hd__buf_4
XFILLER_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _19695_/CLK _18451_/D vssd1 vssd1 vccd1 vccd1 _18451_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ _15663_/A vssd1 vssd1 vccd1 vccd1 _18848_/D sky130_fd_sc_hd__clkbuf_1
X_12875_ _18272_/Q _18271_/Q _18270_/Q _12875_/D vssd1 vssd1 vccd1 vccd1 _12885_/D
+ sky130_fd_sc_hd__and4_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17792__A0 _15149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _16758_/X _19569_/Q _17402_/S vssd1 vssd1 vccd1 vccd1 _17403_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _14519_/A _14613_/X _14603_/X input61/X vssd1 vssd1 vccd1 vccd1 _14615_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15702__S _15708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18382_ _18401_/CLK _18382_/D vssd1 vssd1 vccd1 vccd1 _18382_/Q sky130_fd_sc_hd__dfxtp_1
X_11826_ _11826_/A _11826_/B vssd1 vssd1 vccd1 vccd1 _11826_/Y sky130_fd_sc_hd__nand2_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15594_ _15662_/S vssd1 vssd1 vccd1 vccd1 _15603_/S sky130_fd_sc_hd__buf_2
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _16761_/X _19538_/Q _17341_/S vssd1 vssd1 vccd1 vccd1 _17334_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _14545_/A _14551_/B vssd1 vssd1 vccd1 vccd1 _14545_/Y sky130_fd_sc_hd__nand2_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _12715_/B vssd1 vssd1 vccd1 vccd1 _17762_/S sky130_fd_sc_hd__buf_2
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10708_ _18977_/Q vssd1 vssd1 vccd1 vccd1 _10805_/A sky130_fd_sc_hd__buf_2
X_17264_ _17264_/A vssd1 vssd1 vccd1 vccd1 _19507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14476_ _18509_/Q _19747_/Q _14476_/S vssd1 vssd1 vccd1 vccd1 _14477_/A sky130_fd_sc_hd__mux2_1
X_11688_ _11688_/A _11688_/B _11688_/C _13845_/S vssd1 vssd1 vccd1 vccd1 _13996_/A
+ sky130_fd_sc_hd__and4_2
X_19003_ _19003_/CLK _19003_/D vssd1 vssd1 vccd1 vccd1 _19003_/Q sky130_fd_sc_hd__dfxtp_1
X_16215_ _16283_/S vssd1 vssd1 vccd1 vccd1 _16224_/S sky130_fd_sc_hd__clkbuf_4
X_13427_ _19823_/Q vssd1 vssd1 vccd1 vccd1 _17925_/B sky130_fd_sc_hd__clkbuf_2
X_17195_ _18442_/Q _12559_/X _17201_/S vssd1 vssd1 vccd1 vccd1 _17195_/X sky130_fd_sc_hd__mux2_1
X_10639_ _19509_/Q _19123_/Q _19573_/Q _18729_/Q _10500_/A _09514_/A vssd1 vssd1 vccd1
+ vccd1 _10640_/B sky130_fd_sc_hd__mux4_1
XFILLER_155_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14842__A _14842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09785__B1 _09231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16146_ _16042_/X _19048_/Q _16150_/S vssd1 vssd1 vccd1 vccd1 _16147_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13358_ _19494_/Q _13203_/X _13356_/X _13357_/X vssd1 vssd1 vccd1 vccd1 _13358_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_170_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12309_ _12310_/A _12310_/B vssd1 vssd1 vccd1 vccd1 _12309_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16077_ _16787_/A vssd1 vssd1 vccd1 vccd1 _16077_/X sky130_fd_sc_hd__clkbuf_2
X_13289_ _19870_/Q vssd1 vssd1 vccd1 vccd1 _18247_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__10490__S1 _09587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15028_ _15026_/Y _15027_/X _14969_/A vssd1 vssd1 vccd1 vccd1 _15028_/X sky130_fd_sc_hd__a21o_1
XFILLER_151_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19836_ _19851_/CLK _19836_/D vssd1 vssd1 vccd1 vccd1 _19836_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15086__A1 _11070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_70_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19717_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09671__A _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19767_ _19858_/CLK _19767_/D vssd1 vssd1 vccd1 vccd1 _19767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16979_ _16979_/A vssd1 vssd1 vccd1 vccd1 _19396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14289__A _14289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 io_dbus_rdata[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__11706__A _14431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09520_ _19627_/Q _19465_/Q _18911_/Q _18681_/Q _10389_/S _09483_/X vssd1 vssd1 vccd1
+ vccd1 _09521_/B sky130_fd_sc_hd__mux4_1
XFILLER_65_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18718_ _19725_/CLK _18718_/D vssd1 vssd1 vccd1 vccd1 _18718_/Q sky130_fd_sc_hd__dfxtp_1
X_19698_ _19698_/CLK _19698_/D vssd1 vssd1 vccd1 vccd1 _19698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09451_ _09451_/A vssd1 vssd1 vccd1 vccd1 _09454_/A sky130_fd_sc_hd__buf_2
XANTENNA__10855__C1 _09391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18649_ _19081_/CLK _18649_/D vssd1 vssd1 vccd1 vccd1 _18649_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__14046__C1 _13711_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_85_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19689_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09382_ _10327_/A vssd1 vssd1 vccd1 vccd1 _10144_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18208__B _18214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11441__A _18415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09846__A _09976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_23_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19645_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16510__A1 _15497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10138__A1 _09318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17274__S _17280_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_38_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19725_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_102_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14199__A _14203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09718_ _09712_/A _09715_/X _09717_/X _09708_/X vssd1 vssd1 vccd1 vccd1 _09718_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11616__A _11688_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11638__A1 _18563_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10990_ _10821_/X _10981_/Y _10985_/Y _10989_/Y _09243_/A vssd1 vssd1 vccd1 vccd1
+ _10990_/X sky130_fd_sc_hd__o311a_1
XFILLER_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11335__B _14274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09649_ _09649_/A _09649_/B vssd1 vssd1 vccd1 vccd1 _09649_/X sky130_fd_sc_hd__or2_1
XFILLER_83_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10310__A1 _10313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12660_ _12660_/A vssd1 vssd1 vccd1 vccd1 _13104_/B sky130_fd_sc_hd__buf_2
XFILLER_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _18570_/Q vssd1 vssd1 vccd1 vccd1 _14553_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12591_ _19777_/Q _12590_/X _12628_/A vssd1 vssd1 vccd1 vccd1 _12591_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14330_ _18456_/Q _11460_/A _14319_/Y _14329_/X vssd1 vssd1 vccd1 vccd1 _18456_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11542_ _14999_/A vssd1 vssd1 vccd1 vccd1 _11542_/X sky130_fd_sc_hd__buf_2
XANTENNA__17957__B _19769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15001__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17449__S _17457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11070__B _12462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14261_ _14265_/A _14265_/B vssd1 vssd1 vccd1 vccd1 _14261_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16353__S _16355_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11473_ _11528_/B vssd1 vssd1 vccd1 vccd1 _11474_/B sky130_fd_sc_hd__clkbuf_2
X_16000_ _16000_/A vssd1 vssd1 vccd1 vccd1 _18998_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input70_A io_irq_spi_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ _13121_/X _13202_/Y _13211_/X _13135_/X _18625_/Q vssd1 vssd1 vccd1 vccd1
+ _13212_/X sky130_fd_sc_hd__a32o_4
X_10424_ _10477_/A _10424_/B vssd1 vssd1 vccd1 vccd1 _10424_/X sky130_fd_sc_hd__or2_1
X_14192_ _14192_/A _14192_/B vssd1 vssd1 vccd1 vccd1 _14192_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13143_ _18685_/Q _12671_/X _13141_/X _13142_/X vssd1 vssd1 vccd1 vccd1 _13143_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__13278__A _18632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10355_ _11088_/S vssd1 vssd1 vccd1 vccd1 _11087_/S sky130_fd_sc_hd__buf_2
XFILLER_125_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13315__A1 _12598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17951_ _17954_/B _17954_/C _17950_/X vssd1 vssd1 vccd1 vccd1 _17951_/Y sky130_fd_sc_hd__a21oi_1
X_13074_ _18110_/B _18110_/C _13063_/X vssd1 vssd1 vccd1 vccd1 _13074_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_151_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _09621_/A _10276_/Y _10281_/X _10285_/Y _09393_/A vssd1 vssd1 vccd1 vccd1
+ _10286_/X sky130_fd_sc_hd__o311a_2
XFILLER_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16902_ _19363_/Q _16718_/X _16902_/S vssd1 vssd1 vccd1 vccd1 _16903_/A sky130_fd_sc_hd__mux2_1
X_12025_ _12105_/A vssd1 vssd1 vccd1 vccd1 _12155_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17882_ _17882_/A _17882_/B vssd1 vssd1 vccd1 vccd1 _17883_/A sky130_fd_sc_hd__or2_1
XFILLER_78_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12910__A _18282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09491__A _10500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19621_ _19720_/CLK _19621_/D vssd1 vssd1 vccd1 vccd1 _19621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16833_ _16832_/X _19334_/Q _16839_/S vssd1 vssd1 vccd1 vccd1 _16834_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19552_ _19584_/CLK _19552_/D vssd1 vssd1 vccd1 vccd1 _19552_/Q sky130_fd_sc_hd__dfxtp_1
X_16764_ _16764_/A vssd1 vssd1 vccd1 vccd1 _19312_/D sky130_fd_sc_hd__clkbuf_1
X_13976_ _13984_/A _13984_/B vssd1 vssd1 vccd1 vccd1 _13976_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15715_ _18871_/Q _15561_/X _15719_/S vssd1 vssd1 vccd1 vccd1 _15716_/A sky130_fd_sc_hd__mux2_1
X_18503_ _18506_/CLK _18503_/D vssd1 vssd1 vccd1 vccd1 _18503_/Q sky130_fd_sc_hd__dfxtp_2
X_12927_ _12930_/C _12930_/D _18286_/Q vssd1 vssd1 vccd1 vccd1 _12927_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10837__C1 _09482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19483_ _19682_/CLK _19483_/D vssd1 vssd1 vccd1 vccd1 _19483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16695_ _16695_/A vssd1 vssd1 vccd1 vccd1 _19291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15646_ _15646_/A vssd1 vssd1 vccd1 vccd1 _18840_/D sky130_fd_sc_hd__clkbuf_1
X_18434_ _19695_/CLK _18434_/D vssd1 vssd1 vccd1 vccd1 _18434_/Q sky130_fd_sc_hd__dfxtp_4
X_12858_ _18267_/Q vssd1 vssd1 vccd1 vccd1 _12863_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18365_ _18395_/CLK _18365_/D vssd1 vssd1 vccd1 vccd1 _18365_/Q sky130_fd_sc_hd__dfxtp_1
X_11809_ _11075_/A _18496_/Q _11840_/A vssd1 vssd1 vccd1 vccd1 _11843_/A sky130_fd_sc_hd__mux2_8
XFILLER_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12054__B2 _12483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15577_ _16832_/A vssd1 vssd1 vccd1 vccd1 _15577_/X sky130_fd_sc_hd__clkbuf_2
X_12789_ _15413_/A _12789_/B _12789_/C _12789_/D vssd1 vssd1 vccd1 vccd1 _12790_/D
+ sky130_fd_sc_hd__or4_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _17316_/A vssd1 vssd1 vccd1 vccd1 _19531_/D sky130_fd_sc_hd__clkbuf_1
X_14528_ _14589_/B vssd1 vssd1 vccd1 vccd1 _14582_/B sky130_fd_sc_hd__clkbuf_2
X_18296_ _18298_/CLK _18296_/D vssd1 vssd1 vccd1 vccd1 _18296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17247_ _17391_/B _17535_/B vssd1 vssd1 vccd1 vccd1 _17304_/A sky130_fd_sc_hd__nor2_4
XANTENNA__17359__S _17363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14459_ _18501_/Q _19739_/Q _14465_/S vssd1 vssd1 vccd1 vccd1 _14460_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14572__A _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17178_ _18437_/Q _12713_/X _17184_/S vssd1 vssd1 vccd1 vccd1 _17178_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14751__B1 _14750_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16129_ _16128_/X _19043_/Q _16129_/S vssd1 vssd1 vccd1 vccd1 _16130_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12092__A _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10463__S1 _10368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18245__A1 _18247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19819_ _19822_/CLK _19819_/D vssd1 vssd1 vccd1 vccd1 _19819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14806__A1 _11542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09503_ _09486_/X _09493_/Y _09501_/Y _10227_/A vssd1 vssd1 vccd1 vccd1 _09503_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16438__S _16442_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14747__A _18429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09434_ _09434_/A vssd1 vssd1 vccd1 vccd1 _09434_/X sky130_fd_sc_hd__clkbuf_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09365_ _19274_/Q _19045_/Q _18976_/Q _19370_/Q _09369_/S _09370_/A vssd1 vssd1 vccd1
+ vccd1 _09366_/B sky130_fd_sc_hd__mux4_1
XFILLER_162_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10056__B1 _10068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__A _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09296_ _18574_/Q vssd1 vssd1 vccd1 vccd1 _11516_/A sky130_fd_sc_hd__inv_2
XFILLER_166_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17269__S _17269_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09749__B1 _09621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09576__A _10329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10454__S1 _10245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11110__S _11110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15298__A1 _15181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10140_ _10140_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10140_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_165_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput170 _17862_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[4] sky130_fd_sc_hd__buf_2
X_10071_ _10064_/X _10066_/X _10068_/X _10070_/X _09395_/A vssd1 vssd1 vccd1 vccd1
+ _10071_/X sky130_fd_sc_hd__a221o_1
XFILLER_102_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12730__A _18205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09921__B1 _09231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13830_ _11022_/X _13736_/X _13825_/X _13829_/X vssd1 vssd1 vccd1 vccd1 _18427_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_63_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13761_ _13761_/A vssd1 vssd1 vccd1 vccd1 _13999_/S sky130_fd_sc_hd__clkbuf_2
X_10973_ _10973_/A _10973_/B vssd1 vssd1 vccd1 vccd1 _10973_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18129__A _18173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15500_ _16755_/A vssd1 vssd1 vccd1 vccd1 _15500_/X sky130_fd_sc_hd__buf_2
X_12712_ _12712_/A vssd1 vssd1 vccd1 vccd1 _12712_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16480_ _16103_/X _19200_/Q _16486_/S vssd1 vssd1 vccd1 vccd1 _16481_/A sky130_fd_sc_hd__mux2_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _13684_/X _13691_/X _13991_/S vssd1 vssd1 vccd1 vccd1 _13692_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15431_ _18759_/Q _15159_/X _15437_/S vssd1 vssd1 vccd1 vccd1 _15432_/A sky130_fd_sc_hd__mux2_1
X_12643_ _12643_/A vssd1 vssd1 vccd1 vccd1 _15242_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18150_ _19837_/Q _18150_/B vssd1 vssd1 vccd1 vccd1 _18156_/C sky130_fd_sc_hd__and2_1
XANTENNA__14981__A0 _18449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15362_ _18730_/Q _15168_/X _15362_/S vssd1 vssd1 vccd1 vccd1 _15363_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12574_ _17895_/A vssd1 vssd1 vccd1 vccd1 _12574_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_169_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11795__A0 _11787_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10598__A1 _09529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17101_ _17101_/A vssd1 vssd1 vccd1 vccd1 _19450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14313_ _14310_/B _14308_/B _14003_/X _14311_/X _14312_/X vssd1 vssd1 vccd1 vccd1
+ _14314_/B sky130_fd_sc_hd__o221a_1
X_18081_ _19813_/Q _18077_/B _18080_/Y vssd1 vssd1 vccd1 vccd1 _19813_/D sky130_fd_sc_hd__o21a_1
X_11525_ _13578_/A _12466_/B vssd1 vssd1 vccd1 vccd1 _13587_/A sky130_fd_sc_hd__nor2_2
XANTENNA__15488__A _16430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15293_ _15293_/A vssd1 vssd1 vccd1 vccd1 _18699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10693__S1 _09512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17032_ _19420_/Q _16696_/X _17036_/S vssd1 vssd1 vccd1 vccd1 _17033_/A sky130_fd_sc_hd__mux2_1
X_14244_ _14037_/X _14019_/X _14243_/Y _13737_/A vssd1 vssd1 vccd1 vccd1 _14244_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09486__A _10384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11456_ _14737_/A _14431_/C _14120_/A vssd1 vssd1 vccd1 vccd1 _11457_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10407_ _10438_/A _10406_/X _09411_/A vssd1 vssd1 vccd1 vccd1 _10407_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_171_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14175_ _18443_/Q _13736_/X _14163_/Y _14174_/X vssd1 vssd1 vccd1 vccd1 _18443_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_125_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16811__S _16823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11387_ _18422_/Q vssd1 vssd1 vccd1 vccd1 _14802_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_125_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15289__A1 _15168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13126_ _13270_/B vssd1 vssd1 vccd1 vccd1 _13126_/X sky130_fd_sc_hd__clkbuf_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10338_ _19644_/Q _19061_/Q _19098_/Q _18704_/Q _11188_/S _09610_/A vssd1 vssd1 vccd1
+ vccd1 _10338_/X sky130_fd_sc_hd__mux4_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ _19597_/CLK _18983_/D vssd1 vssd1 vccd1 vccd1 _18983_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13736__A _14120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17934_ _19763_/Q _17934_/B _17934_/C vssd1 vssd1 vccd1 vccd1 _17935_/C sky130_fd_sc_hd__and3_1
X_13057_ _17999_/A vssd1 vssd1 vccd1 vccd1 _17948_/A sky130_fd_sc_hd__clkbuf_2
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10269_ _19613_/Q _19451_/Q _18897_/Q _18667_/Q _09794_/A _09145_/A vssd1 vssd1 vccd1
+ vccd1 _10270_/B sky130_fd_sc_hd__mux4_1
XANTENNA__16112__A _16822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12008_ _12008_/A _12008_/B vssd1 vssd1 vccd1 vccd1 _12010_/A sky130_fd_sc_hd__xor2_4
XFILLER_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17865_ _18225_/A vssd1 vssd1 vccd1 vccd1 _17874_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_66_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19604_ _19636_/CLK _19604_/D vssd1 vssd1 vccd1 vccd1 _19604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16816_ _16816_/A vssd1 vssd1 vccd1 vccd1 _16816_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17796_ _17853_/S vssd1 vssd1 vccd1 vccd1 _17805_/S sky130_fd_sc_hd__buf_2
XFILLER_47_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19535_ _19537_/CLK _19535_/D vssd1 vssd1 vccd1 vccd1 _19535_/Q sky130_fd_sc_hd__dfxtp_1
X_13959_ _13810_/A _13953_/X _13958_/X vssd1 vssd1 vccd1 vccd1 _13959_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_34_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16747_ _16743_/X _19307_/Q _16759_/S vssd1 vssd1 vccd1 vccd1 _16748_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11406__D _11406_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18039__A _18170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19466_ _19660_/CLK _19466_/D vssd1 vssd1 vccd1 vccd1 _19466_/Q sky130_fd_sc_hd__dfxtp_1
X_16678_ _19286_/Q _16677_/X _16687_/S vssd1 vssd1 vccd1 vccd1 _16679_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18417_ _18509_/CLK _18417_/D vssd1 vssd1 vccd1 vccd1 _18417_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__17878__A _17878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12027__B2 _12482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15629_ _15629_/A vssd1 vssd1 vccd1 vccd1 _18832_/D sky130_fd_sc_hd__clkbuf_1
X_19397_ _19397_/CLK _19397_/D vssd1 vssd1 vccd1 vccd1 _19397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09150_ _19691_/Q vssd1 vssd1 vccd1 vccd1 _11028_/S sky130_fd_sc_hd__buf_2
X_18348_ _18386_/CLK _18348_/D vssd1 vssd1 vccd1 vccd1 _18348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17089__S _17097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18279_ _18298_/CLK _18279_/D vssd1 vssd1 vccd1 vccd1 _18279_/Q sky130_fd_sc_hd__dfxtp_1
X_09081_ _18557_/Q _18556_/Q _18555_/Q _18554_/Q vssd1 vssd1 vccd1 vccd1 _09088_/A
+ sky130_fd_sc_hd__or4bb_1
XANTENNA__10684__S1 _09139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput50 io_ibus_inst[24] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_2
XFILLER_147_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput61 io_ibus_inst[5] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_1
Xinput72 reset vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__buf_4
XFILLER_156_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09983_ _10200_/S vssd1 vssd1 vccd1 vccd1 _09983_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15337__S _15337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12550__A _12628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11166__A _11166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12266__A1 _12246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11069__A2 _12460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16168__S _16172_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09417_ _09421_/A _09417_/B vssd1 vssd1 vccd1 vccd1 _09417_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_91_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15800__S _15802_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09348_ _09928_/A vssd1 vssd1 vccd1 vccd1 _09367_/S sky130_fd_sc_hd__buf_2
XANTENNA__11777__B1 _11970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09279_ _11046_/B vssd1 vssd1 vccd1 vccd1 _09280_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13518__A1 _18415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11310_ _11475_/A _11585_/B _11495_/B vssd1 vssd1 vccd1 vccd1 _11310_/X sky130_fd_sc_hd__or3_1
XANTENNA__13518__B2 _14431_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12290_ _12371_/A _12290_/B vssd1 vssd1 vccd1 vccd1 _12290_/X sky130_fd_sc_hd__xor2_4
XFILLER_153_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11241_ _11239_/Y _11135_/X _10413_/A _11263_/A vssd1 vssd1 vccd1 vccd1 _11266_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10245__A _10245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11172_ _11166_/A _11169_/X _11171_/X _09708_/X vssd1 vssd1 vccd1 vccd1 _11172_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10123_ _10007_/X _10118_/X _10120_/X _10122_/X _09135_/A vssd1 vssd1 vccd1 vccd1
+ _10123_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15980_ _15980_/A vssd1 vssd1 vccd1 vccd1 _18989_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09753__B _12500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12460__A _12460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13151__C1 _13102_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10054_ _09880_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _10054_/X sky130_fd_sc_hd__and2b_1
X_14931_ _14931_/A vssd1 vssd1 vccd1 vccd1 _18604_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input33_A io_dbus_valid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17650_ _17645_/A _17649_/C _14366_/X vssd1 vssd1 vccd1 vccd1 _17651_/B sky130_fd_sc_hd__o21ai_1
X_14862_ _17662_/A _14861_/A _14840_/B _18471_/Q vssd1 vssd1 vccd1 vccd1 _14863_/C
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11507__C _13529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13813_ _13968_/S _13818_/B vssd1 vssd1 vccd1 vccd1 _13813_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16601_ _19256_/Q vssd1 vssd1 vccd1 vccd1 _16602_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_75_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17581_ _17592_/A vssd1 vssd1 vccd1 vccd1 _17590_/S sky130_fd_sc_hd__buf_4
XANTENNA__16078__S _16081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14793_ _14792_/X _18593_/Q _14822_/S vssd1 vssd1 vccd1 vccd1 _14794_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16532_ _19223_/Q _15529_/X _16536_/S vssd1 vssd1 vccd1 vccd1 _16533_/A sky130_fd_sc_hd__mux2_1
X_19320_ _19610_/CLK _19320_/D vssd1 vssd1 vccd1 vccd1 _19320_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10268__B1 _09214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13744_ _13993_/A vssd1 vssd1 vccd1 vccd1 _13881_/S sky130_fd_sc_hd__clkbuf_2
X_10956_ _10956_/A _10956_/B vssd1 vssd1 vccd1 vccd1 _10956_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16463_ _16463_/A vssd1 vssd1 vccd1 vccd1 _19192_/D sky130_fd_sc_hd__clkbuf_1
X_19251_ _19659_/CLK _19251_/D vssd1 vssd1 vccd1 vccd1 _19251_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12009__A1 _18503_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13675_ _13669_/X _13673_/X _13877_/S vssd1 vssd1 vccd1 vccd1 _13675_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10887_ _10887_/A _10887_/B vssd1 vssd1 vccd1 vccd1 _10887_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18202_ _19854_/Q _18200_/B _18201_/Y vssd1 vssd1 vccd1 vccd1 _19854_/D sky130_fd_sc_hd__o21a_1
XFILLER_148_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15414_ _16992_/A vssd1 vssd1 vccd1 vccd1 _17535_/B sky130_fd_sc_hd__clkbuf_4
X_12626_ _19678_/Q _12703_/A _12742_/A _18402_/Q _12625_/X vssd1 vssd1 vccd1 vccd1
+ _12626_/X sky130_fd_sc_hd__a221o_1
X_19182_ _19632_/CLK _19182_/D vssd1 vssd1 vccd1 vccd1 _19182_/Q sky130_fd_sc_hd__dfxtp_1
X_16394_ _19162_/Q _15538_/X _16402_/S vssd1 vssd1 vccd1 vccd1 _16395_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18133_ _19831_/Q _19830_/Q _19829_/Q _18133_/D vssd1 vssd1 vccd1 vccd1 _18142_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_12_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15345_ _18722_/Q _15143_/X _15351_/S vssd1 vssd1 vccd1 vccd1 _15346_/A sky130_fd_sc_hd__mux2_1
X_12557_ _12557_/A vssd1 vssd1 vccd1 vccd1 _12712_/A sky130_fd_sc_hd__buf_2
XFILLER_8_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18064_ _19807_/Q _18061_/B _18063_/Y vssd1 vssd1 vccd1 vccd1 _19807_/D sky130_fd_sc_hd__o21a_1
XFILLER_8_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11508_ _13521_/B _14089_/A _11508_/C vssd1 vssd1 vccd1 vccd1 _11522_/B sky130_fd_sc_hd__and3_1
XFILLER_145_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15276_ _18692_/Q _15149_/X _15278_/S vssd1 vssd1 vccd1 vccd1 _15277_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12488_ _12488_/A _12497_/B vssd1 vssd1 vccd1 vccd1 _12488_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09189__A1 _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17015_ _17015_/A vssd1 vssd1 vccd1 vccd1 _19412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14227_ _14227_/A _14227_/B vssd1 vssd1 vccd1 vccd1 _14227_/Y sky130_fd_sc_hd__nand2_1
X_11439_ _18418_/Q _18417_/Q _18419_/Q vssd1 vssd1 vccd1 vccd1 _12688_/C sky130_fd_sc_hd__or3b_1
XFILLER_160_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16541__S _16547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14158_ _14150_/X _14137_/Y _14157_/X vssd1 vssd1 vccd1 vccd1 _14158_/X sky130_fd_sc_hd__a21o_1
XFILLER_152_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _15242_/A _13536_/A _13442_/D vssd1 vssd1 vccd1 vccd1 _13109_/X sky130_fd_sc_hd__and3_2
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18966_ _19717_/CLK _18966_/D vssd1 vssd1 vccd1 vccd1 _18966_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ _14089_/A _14089_/B vssd1 vssd1 vccd1 vccd1 _14089_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15682__A1 _15513_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17917_ _19805_/Q _19807_/Q _19806_/Q _18054_/A vssd1 vssd1 vccd1 vccd1 _18062_/A
+ sky130_fd_sc_hd__and4_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11379__B1_N _09624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18897_ _19581_/CLK _18897_/D vssd1 vssd1 vccd1 vccd1 _18897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17372__S _17374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17848_ _17848_/A vssd1 vssd1 vccd1 vccd1 _19724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11417__C _11821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17779_ _17779_/A _17779_/B vssd1 vssd1 vccd1 vccd1 _17780_/A sky130_fd_sc_hd__and2_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19518_ _19613_/CLK _19518_/D vssd1 vssd1 vccd1 vccd1 _19518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_113_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19449_ _19609_/CLK _19449_/D vssd1 vssd1 vccd1 vccd1 _19449_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16716__S _16719_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09202_ _10212_/A vssd1 vssd1 vccd1 vccd1 _10074_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ _09133_/A vssd1 vssd1 vccd1 vccd1 _09134_/A sky130_fd_sc_hd__buf_4
XFILLER_120_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09854__A _09854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15067__S _15077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _19651_/Q _19068_/Q _19105_/Q _18711_/Q _09803_/A _09936_/X vssd1 vssd1 vccd1
+ vccd1 _09966_/X sky130_fd_sc_hd__mux4_1
XANTENNA__15673__A1 _15500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _09898_/A _12499_/A vssd1 vssd1 vccd1 vccd1 _11151_/A sky130_fd_sc_hd__nand2_1
XFILLER_134_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _18430_/Q vssd1 vssd1 vccd1 vccd1 _10810_/X sky130_fd_sc_hd__buf_6
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _11790_/A vssd1 vssd1 vccd1 vccd1 _11790_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17178__A1 _12713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10741_ _09629_/A _10736_/Y _10738_/Y _10740_/X vssd1 vssd1 vccd1 vccd1 _10741_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10896__S1 _10726_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15530__S _15536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13460_ _18390_/Q _13110_/A _13464_/S vssd1 vssd1 vccd1 vccd1 _13461_/A sky130_fd_sc_hd__mux2_1
X_10672_ _19250_/Q _19021_/Q _18952_/Q _19346_/Q _10614_/X _10616_/X vssd1 vssd1 vccd1
+ vccd1 _10672_/X sky130_fd_sc_hd__mux4_2
X_12411_ _12434_/B _12411_/B _12411_/C vssd1 vssd1 vccd1 vccd1 _12411_/X sky130_fd_sc_hd__and3b_1
XFILLER_138_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13391_ _18295_/Q _13126_/X _13127_/X _18378_/Q vssd1 vssd1 vccd1 vccd1 _13391_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15130_ hold3/A _13873_/X _15125_/X _11200_/A vssd1 vssd1 vccd1 vccd1 _18648_/D sky130_fd_sc_hd__a22o_1
X_12342_ _12193_/X _12340_/Y _12393_/C _12186_/A vssd1 vssd1 vccd1 vccd1 _12342_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_138_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15061_ _14958_/A _13422_/B _15060_/X _14893_/A vssd1 vssd1 vccd1 vccd1 _15061_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17457__S _17457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12273_ _17611_/B vssd1 vssd1 vccd1 vccd1 _17693_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__16361__S _16369_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18142__A _19834_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12175__B1 _12057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14012_ _14115_/A vssd1 vssd1 vccd1 vccd1 _14012_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13911__A1 _11704_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ _11224_/A vssd1 vssd1 vccd1 vccd1 _11224_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18820_ _19691_/CLK _18820_/D vssd1 vssd1 vccd1 vccd1 _18820_/Q sky130_fd_sc_hd__dfxtp_1
X_11155_ _11168_/A _11155_/B vssd1 vssd1 vccd1 vccd1 _11155_/X sky130_fd_sc_hd__or2_1
XFILLER_68_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13717__C _13720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10106_ _19648_/Q _19065_/Q _19102_/Q _18708_/Q _10094_/X _10103_/X vssd1 vssd1 vccd1
+ vccd1 _10107_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18751_ _19713_/CLK _18751_/D vssd1 vssd1 vccd1 vccd1 _18751_/Q sky130_fd_sc_hd__dfxtp_1
X_15963_ _16031_/S vssd1 vssd1 vccd1 vccd1 _15972_/S sky130_fd_sc_hd__clkbuf_4
X_11086_ _11097_/A _11086_/B vssd1 vssd1 vccd1 vccd1 _11086_/X sky130_fd_sc_hd__or2_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17702_ _17701_/A _17701_/C _17701_/B vssd1 vssd1 vccd1 vccd1 _17703_/B sky130_fd_sc_hd__o21ai_1
X_10037_ _10042_/A _10037_/B vssd1 vssd1 vccd1 vccd1 _10037_/X sky130_fd_sc_hd__or2_1
XFILLER_64_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14914_ _14969_/A _14911_/X _14932_/C _14913_/Y vssd1 vssd1 vccd1 vccd1 _14914_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_49_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15894_ _14772_/X _18950_/Q _15902_/S vssd1 vssd1 vccd1 vccd1 _15895_/A sky130_fd_sc_hd__mux2_1
X_18682_ _19647_/CLK _18682_/D vssd1 vssd1 vccd1 vccd1 _18682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17633_ _17632_/A _17632_/C _14786_/A vssd1 vssd1 vccd1 vccd1 _17634_/B sky130_fd_sc_hd__o21ai_1
X_14845_ _14845_/A _14845_/B vssd1 vssd1 vccd1 vccd1 _16677_/A sky130_fd_sc_hd__nor2_8
XFILLER_84_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17564_ _19641_/Q _16784_/A _17568_/S vssd1 vssd1 vccd1 vccd1 _17565_/A sky130_fd_sc_hd__mux2_1
X_14776_ _14786_/A _14786_/C vssd1 vssd1 vccd1 vccd1 _14776_/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11988_ _12412_/B vssd1 vssd1 vccd1 vccd1 _12098_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10336__S0 _10125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19303_ _19626_/CLK _19303_/D vssd1 vssd1 vccd1 vccd1 _19303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16515_ _16515_/A vssd1 vssd1 vccd1 vccd1 _19215_/D sky130_fd_sc_hd__clkbuf_1
X_13727_ _14150_/A _13706_/Y _13723_/X _13726_/X vssd1 vssd1 vccd1 vccd1 _13727_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_90_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10939_ _11056_/A vssd1 vssd1 vccd1 vccd1 _11060_/A sky130_fd_sc_hd__clkbuf_1
X_17495_ _17495_/A vssd1 vssd1 vccd1 vccd1 _19610_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15440__S _15448_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19234_ _19557_/CLK _19234_/D vssd1 vssd1 vccd1 vccd1 _19234_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17221__A _17221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13658_ _13658_/A vssd1 vssd1 vccd1 vccd1 _13658_/X sky130_fd_sc_hd__clkbuf_2
X_16446_ _16446_/A vssd1 vssd1 vccd1 vccd1 _19184_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12609_ _19487_/Q _12669_/A _12674_/A _18401_/Q _12608_/X vssd1 vssd1 vccd1 vccd1
+ _12609_/X sky130_fd_sc_hd__a221o_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16377_ _16377_/A vssd1 vssd1 vccd1 vccd1 _19154_/D sky130_fd_sc_hd__clkbuf_1
X_19165_ _19165_/CLK _19165_/D vssd1 vssd1 vccd1 vccd1 _19165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10639__S1 _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13589_ _14332_/B _13729_/B vssd1 vssd1 vccd1 vccd1 _13589_/X sky130_fd_sc_hd__xor2_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18116_ _18119_/B _18119_/C _18082_/X vssd1 vssd1 vccd1 vccd1 _18116_/Y sky130_fd_sc_hd__a21oi_1
X_15328_ _15328_/A vssd1 vssd1 vccd1 vccd1 _18715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19096_ _19546_/CLK _19096_/D vssd1 vssd1 vccd1 vccd1 _19096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12084__B _13604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15259_ _15258_/X _17149_/B _11822_/X vssd1 vssd1 vccd1 vccd1 _15259_/Y sky130_fd_sc_hd__o21ai_1
X_18047_ _18071_/A _18051_/C vssd1 vssd1 vccd1 vccd1 _18047_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16271__S _16279_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14580__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09820_ _18873_/Q _19331_/Q _09955_/A vssd1 vssd1 vccd1 vccd1 _09821_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13196__A _18624_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09751_ _18452_/Q vssd1 vssd1 vccd1 vccd1 _09751_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13666__A0 _12401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18949_ _19700_/CLK _18949_/D vssd1 vssd1 vccd1 vccd1 _18949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09682_ _11123_/A _09680_/X _09681_/X vssd1 vssd1 vccd1 vccd1 _09682_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10575__S0 _11088_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13418__A0 _11406_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17830__S _17838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10194__A1_N _18444_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09116_ _11343_/B vssd1 vssd1 vccd1 vccd1 _11361_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16181__S _16183_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09584__A _10328_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10707__A1 _10887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09573__A1 _09214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10802__S1 _10772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09949_ _09415_/X _09942_/X _09944_/X _09948_/X _09395_/X vssd1 vssd1 vccd1 vccd1
+ _09949_/X sky130_fd_sc_hd__a311o_4
XANTENNA__13657__A0 _14265_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12960_ _18297_/Q _12959_/B _12574_/X vssd1 vssd1 vccd1 vccd1 _12961_/B sky130_fd_sc_hd__o21ai_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ _14587_/A _12173_/A _11911_/C vssd1 vssd1 vccd1 vccd1 _11911_/X sky130_fd_sc_hd__and3_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12891_ _12895_/C _12893_/C _12890_/Y vssd1 vssd1 vccd1 vccd1 _18276_/D sky130_fd_sc_hd__o21a_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _18564_/Q _14613_/X _14622_/X input35/X vssd1 vssd1 vccd1 vccd1 _14631_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11354__A _11513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _11842_/A _13658_/A vssd1 vssd1 vccd1 vccd1 _11846_/A sky130_fd_sc_hd__xor2_4
XANTENNA__10891__B1 _10793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10318__S0 _09701_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _18541_/Q _14550_/X _14559_/X _14560_/X vssd1 vssd1 vccd1 vccd1 _18541_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11773_ _11966_/B _15095_/B vssd1 vssd1 vccd1 vccd1 _11911_/C sky130_fd_sc_hd__nor2_2
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _18414_/Q _13437_/Y _13512_/S vssd1 vssd1 vccd1 vccd1 _13513_/A sky130_fd_sc_hd__mux2_1
X_16300_ _16300_/A vssd1 vssd1 vccd1 vccd1 _19120_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09759__A _10076_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10724_ _10724_/A vssd1 vssd1 vccd1 vccd1 _10724_/X sky130_fd_sc_hd__buf_4
X_17280_ _19515_/Q _16686_/X _17280_/S vssd1 vssd1 vccd1 vccd1 _17281_/A sky130_fd_sc_hd__mux2_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _18516_/Q _19754_/Q _14498_/S vssd1 vssd1 vccd1 vccd1 _14493_/A sky130_fd_sc_hd__mux2_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17571__A1 _16793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16231_ _16058_/X _19090_/Q _16235_/S vssd1 vssd1 vccd1 vccd1 _16232_/A sky130_fd_sc_hd__mux2_1
X_13443_ _13499_/A vssd1 vssd1 vccd1 vccd1 _13512_/S sky130_fd_sc_hd__clkbuf_2
X_10655_ _10762_/A _10654_/X _09517_/A vssd1 vssd1 vccd1 vccd1 _10655_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16162_ _16162_/A vssd1 vssd1 vccd1 vccd1 _19055_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13374_ _19495_/Q _13203_/X _13369_/X _13370_/X _13373_/X vssd1 vssd1 vccd1 vccd1
+ _15018_/B sky130_fd_sc_hd__a2111o_2
XFILLER_139_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10586_ _18762_/Q _18991_/Q _18922_/Q _19220_/Q _10500_/A _09514_/A vssd1 vssd1 vccd1
+ vccd1 _10587_/B sky130_fd_sc_hd__mux4_1
XFILLER_10_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15113_ _18635_/Q _15109_/X _15111_/X _10299_/A vssd1 vssd1 vccd1 vccd1 _18635_/D
+ sky130_fd_sc_hd__a22o_1
X_12325_ _12419_/A _12325_/B vssd1 vssd1 vccd1 vccd1 _14274_/B sky130_fd_sc_hd__nand2_4
XFILLER_154_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16091__S _16097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16093_ _16803_/A vssd1 vssd1 vccd1 vccd1 _16093_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09239__S1 _09149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15044_ _16835_/A vssd1 vssd1 vccd1 vccd1 _15044_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09494__A _18977_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12256_ _12256_/A vssd1 vssd1 vccd1 vccd1 _14241_/A sky130_fd_sc_hd__buf_2
XFILLER_141_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12632__B _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11529__A _12505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11207_ _11207_/A vssd1 vssd1 vccd1 vccd1 _11284_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09564__A1 _09214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19852_ _19871_/CLK _19852_/D vssd1 vssd1 vccd1 vccd1 _19852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12187_ _19747_/Q _12215_/C vssd1 vssd1 vccd1 vccd1 _12188_/B sky130_fd_sc_hd__nand2_1
XFILLER_122_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18803_ _19551_/CLK _18803_/D vssd1 vssd1 vccd1 vccd1 _18803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11138_ _11235_/A _11239_/A _11235_/C _10300_/A _11137_/X vssd1 vssd1 vccd1 vccd1
+ _11230_/C sky130_fd_sc_hd__a311o_1
X_19783_ _19790_/CLK _19783_/D vssd1 vssd1 vccd1 vccd1 _19783_/Q sky130_fd_sc_hd__dfxtp_1
X_16995_ _19403_/Q _16639_/X _17003_/S vssd1 vssd1 vccd1 vccd1 _16996_/A sky130_fd_sc_hd__mux2_1
X_18734_ _19546_/CLK _18734_/D vssd1 vssd1 vccd1 vccd1 _18734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11069_ _11619_/A _12460_/A _11047_/X _12458_/A vssd1 vssd1 vccd1 vccd1 _11257_/A
+ sky130_fd_sc_hd__a22o_1
X_15946_ _15055_/X _18974_/Q _15946_/S vssd1 vssd1 vccd1 vccd1 _15947_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18665_ _19609_/CLK _18665_/D vssd1 vssd1 vccd1 vccd1 _18665_/Q sky130_fd_sc_hd__dfxtp_1
X_15877_ _15877_/A vssd1 vssd1 vccd1 vccd1 _18943_/D sky130_fd_sc_hd__clkbuf_1
X_17616_ _17616_/A vssd1 vssd1 vccd1 vccd1 _19661_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14828_ _17645_/A _14366_/X _14796_/B _18468_/Q vssd1 vssd1 vccd1 vccd1 _14829_/C
+ sky130_fd_sc_hd__a31o_1
X_18596_ _19285_/CLK _18596_/D vssd1 vssd1 vccd1 vccd1 _18596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17547_ _17547_/A vssd1 vssd1 vccd1 vccd1 _19633_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16266__S _16268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14575__A _14575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14759_ input27/X _14703_/X _14758_/X _14732_/X vssd1 vssd1 vccd1 vccd1 _16654_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17478_ _17478_/A vssd1 vssd1 vccd1 vccd1 _19602_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19217_ _19539_/CLK _19217_/D vssd1 vssd1 vccd1 vccd1 _19217_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14376__A1 _18502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16429_ _16429_/A vssd1 vssd1 vccd1 vccd1 _19178_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12095__A _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16790__A _16790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19148_ _19598_/CLK _19148_/D vssd1 vssd1 vccd1 vccd1 _19148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17097__S _17097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19079_ _19079_/CLK _19079_/D vssd1 vssd1 vccd1 vccd1 _19079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13336__C1 _13317_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17078__A0 _16761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13351__A2 _13139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17825__S _17827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09803_ _09803_/A vssd1 vssd1 vccd1 vccd1 _09803_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_113_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10796__S0 _10934_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15345__S _15351_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13103__A2 _12731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _09734_/A vssd1 vssd1 vccd1 vccd1 _09734_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09665_ _19528_/Q _19142_/Q _19592_/Q _18748_/Q _10328_/S _10280_/A vssd1 vssd1 vccd1
+ vccd1 _09666_/B sky130_fd_sc_hd__mux4_1
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10322__C1 _09133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17560__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09596_ _10400_/A vssd1 vssd1 vccd1 vccd1 _09671_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10720__S0 _10719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17796__A _17853_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10440_ _10447_/A _10440_/B vssd1 vssd1 vccd1 vccd1 _10440_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10371_ _10477_/A _10371_/B vssd1 vssd1 vccd1 vccd1 _10371_/X sky130_fd_sc_hd__or2_1
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13327__C1 _13326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12110_ _12111_/A _13608_/A vssd1 vssd1 vccd1 vccd1 _12112_/A sky130_fd_sc_hd__and2_1
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13090_ _18341_/Q _13089_/X _13090_/S vssd1 vssd1 vccd1 vccd1 _13091_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17069__A0 _16749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12041_ _12041_/A vssd1 vssd1 vccd1 vccd1 _12041_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_172_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10253__A _11137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15800_ _15044_/X _18909_/Q _15802_/S vssd1 vssd1 vccd1 vccd1 _15801_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16780_ _16780_/A vssd1 vssd1 vccd1 vccd1 _19317_/D sky130_fd_sc_hd__clkbuf_1
X_13992_ _13992_/A vssd1 vssd1 vccd1 vccd1 _13992_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11105__B2 _18439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12943_ _12943_/A _12943_/B _12945_/B vssd1 vssd1 vccd1 vccd1 _18291_/D sky130_fd_sc_hd__nor3_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15731_ _15731_/A vssd1 vssd1 vccd1 vccd1 _18878_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17241__A0 _18456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17470__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18450_ _18632_/CLK _18450_/D vssd1 vssd1 vccd1 vccd1 _18450_/Q sky130_fd_sc_hd__dfxtp_4
X_12874_ _12904_/A _12874_/B _12874_/C vssd1 vssd1 vccd1 vccd1 _18271_/D sky130_fd_sc_hd__nor3_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _18848_/Q _15589_/X _15662_/S vssd1 vssd1 vccd1 vccd1 _15663_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _17401_/A vssd1 vssd1 vccd1 vccd1 _19568_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11825_ _11826_/A _11826_/B vssd1 vssd1 vccd1 vccd1 _11825_/X sky130_fd_sc_hd__or2_1
X_14613_ _14648_/A vssd1 vssd1 vccd1 vccd1 _14613_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18381_ _18381_/CLK _18381_/D vssd1 vssd1 vccd1 vccd1 _18381_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15593_ _15649_/A vssd1 vssd1 vccd1 vccd1 _15662_/S sky130_fd_sc_hd__clkbuf_16
XANTENNA_output102_A _11846_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_7_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12908__A _12997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14544_ _18534_/Q _14522_/X _14543_/Y _14535_/X vssd1 vssd1 vccd1 vccd1 _18534_/D
+ sky130_fd_sc_hd__o211a_1
X_17332_ _17389_/S vssd1 vssd1 vccd1 vccd1 _17341_/S sky130_fd_sc_hd__buf_2
XANTENNA__09489__A _10770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _11563_/X _11751_/X _11754_/X _11755_/Y vssd1 vssd1 vccd1 vccd1 _11756_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_14_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10707_ _10887_/A _10706_/X _10791_/A vssd1 vssd1 vccd1 vccd1 _10707_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17263_ _19507_/Q _16661_/X _17269_/S vssd1 vssd1 vccd1 vccd1 _17264_/A sky130_fd_sc_hd__mux2_1
X_14475_ _14475_/A vssd1 vssd1 vccd1 vccd1 _18508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16814__S _16823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11687_ _12462_/A _11638_/Y _11835_/S vssd1 vssd1 vccd1 vccd1 _13845_/S sky130_fd_sc_hd__mux2_4
X_19002_ _19326_/CLK _19002_/D vssd1 vssd1 vccd1 vccd1 _19002_/Q sky130_fd_sc_hd__dfxtp_1
X_13426_ _13426_/A _18650_/Q vssd1 vssd1 vccd1 vccd1 _13426_/Y sky130_fd_sc_hd__nand2_1
X_16214_ _16270_/A vssd1 vssd1 vccd1 vccd1 _16283_/S sky130_fd_sc_hd__buf_6
X_17194_ _17194_/A vssd1 vssd1 vccd1 vccd1 _19484_/D sky130_fd_sc_hd__clkbuf_1
X_10638_ _10638_/A _10638_/B vssd1 vssd1 vccd1 vccd1 _10638_/Y sky130_fd_sc_hd__nor2_1
XFILLER_167_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16145_ _16145_/A vssd1 vssd1 vccd1 vccd1 _19047_/D sky130_fd_sc_hd__clkbuf_1
X_13357_ _19684_/Q _13251_/X _12743_/X _18408_/Q vssd1 vssd1 vccd1 vccd1 _13357_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13739__A _13845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10569_ _19510_/Q _19124_/Q _19574_/Q _18730_/Q _10466_/S _10559_/A vssd1 vssd1 vccd1
+ vccd1 _10570_/B sky130_fd_sc_hd__mux4_1
XFILLER_170_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13318__C1 _13317_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_4_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19337_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12308_ _14265_/B vssd1 vssd1 vccd1 vccd1 _12310_/B sky130_fd_sc_hd__inv_2
XFILLER_170_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16076_ _16076_/A vssd1 vssd1 vccd1 vccd1 _19026_/D sky130_fd_sc_hd__clkbuf_1
X_13288_ _13288_/A _13288_/B vssd1 vssd1 vccd1 vccd1 _14873_/B sky130_fd_sc_hd__or2_1
XFILLER_108_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15027_ _15027_/A _15037_/C vssd1 vssd1 vccd1 vccd1 _15027_/X sky130_fd_sc_hd__or2_1
XANTENNA__14530__A1 _18562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12239_ _12240_/A _12240_/B vssd1 vssd1 vccd1 vccd1 _12241_/A sky130_fd_sc_hd__nand2_1
XFILLER_130_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19835_ _19838_/CLK _19835_/D vssd1 vssd1 vccd1 vccd1 _19835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19766_ _19858_/CLK _19766_/D vssd1 vssd1 vccd1 vccd1 _19766_/Q sky130_fd_sc_hd__dfxtp_1
X_16978_ _16825_/X _19396_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16979_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14294__B1 _15123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14289__B _14289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput4 io_dbus_rdata[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_2
X_18717_ _19271_/CLK _18717_/D vssd1 vssd1 vccd1 vccd1 _18717_/Q sky130_fd_sc_hd__dfxtp_1
X_15929_ _14964_/X _18966_/Q _15935_/S vssd1 vssd1 vccd1 vccd1 _15930_/A sky130_fd_sc_hd__mux2_1
X_19697_ _19697_/CLK _19697_/D vssd1 vssd1 vccd1 vccd1 _19697_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17232__A0 _18453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09450_ _18879_/Q _19337_/Q _10348_/S vssd1 vssd1 vccd1 vccd1 _09450_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18648_ _19727_/CLK _18648_/D vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_2
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09381_ _09661_/A vssd1 vssd1 vccd1 vccd1 _10327_/A sky130_fd_sc_hd__buf_2
XFILLER_52_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18579_ _18585_/CLK _18579_/D vssd1 vssd1 vccd1 vccd1 _18579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11722__A _11821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12537__B _12537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10702__S0 _10770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10083__A1 _10093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11441__B _18427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09776__A1 _09861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09717_ _10262_/A _09717_/B vssd1 vssd1 vccd1 vccd1 _09717_/X sky130_fd_sc_hd__or2_1
XFILLER_28_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09648_ _19528_/Q _19142_/Q _19592_/Q _18748_/Q _11153_/A _09636_/X vssd1 vssd1 vccd1
+ vccd1 _09649_/B sky130_fd_sc_hd__mux4_1
XFILLER_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09579_ _09661_/A vssd1 vssd1 vccd1 vccd1 _10175_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_161_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11632__A _11688_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11610_ _11610_/A vssd1 vssd1 vccd1 vccd1 _11835_/S sky130_fd_sc_hd__buf_2
XFILLER_35_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _18339_/Q _12531_/Y _12586_/X _12589_/X vssd1 vssd1 vccd1 vccd1 _12590_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11541_ _19080_/Q vssd1 vssd1 vccd1 vccd1 _14999_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14260_ _14260_/A vssd1 vssd1 vccd1 vccd1 _18450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ _11472_/A vssd1 vssd1 vccd1 vccd1 _11474_/A sky130_fd_sc_hd__clkbuf_2
X_13211_ _18625_/Q _13211_/B vssd1 vssd1 vccd1 vccd1 _13211_/X sky130_fd_sc_hd__or2_1
XFILLER_137_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10423_ _18765_/Q _18994_/Q _18925_/Q _19223_/Q _11088_/S _10559_/A vssd1 vssd1 vccd1
+ vccd1 _10424_/B sky130_fd_sc_hd__mux4_1
XFILLER_137_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14191_ _13975_/X _14188_/Y _14190_/X _13982_/X vssd1 vssd1 vccd1 vccd1 _14191_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_125_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12463__A _12463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13142_ _18268_/Q _13126_/X _13127_/A _18351_/Q vssd1 vssd1 vccd1 vccd1 _13142_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input63_A io_ibus_inst[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ _10558_/S vssd1 vssd1 vccd1 vccd1 _11088_/S sky130_fd_sc_hd__buf_6
XFILLER_151_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09519__A1 _09315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13073_ _18334_/Q vssd1 vssd1 vccd1 vccd1 _18110_/B sky130_fd_sc_hd__clkbuf_2
X_17950_ _17993_/A vssd1 vssd1 vccd1 vccd1 _17950_/X sky130_fd_sc_hd__clkbuf_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10285_ _09671_/A _10282_/X _10284_/X vssd1 vssd1 vccd1 vccd1 _10285_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18150__A _19837_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16901_ _16901_/A vssd1 vssd1 vccd1 vccd1 _19362_/D sky130_fd_sc_hd__clkbuf_1
X_12024_ _12024_/A _12323_/A vssd1 vssd1 vccd1 vccd1 _12105_/A sky130_fd_sc_hd__or2_2
XFILLER_78_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_86_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17881_ _17881_/A vssd1 vssd1 vccd1 vccd1 _19741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12910__B _18281_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19620_ _19620_/CLK _19620_/D vssd1 vssd1 vccd1 vccd1 _19620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16832_ _16832_/A vssd1 vssd1 vccd1 vccd1 _16832_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10711__A _10711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19551_ _19551_/CLK _19551_/D vssd1 vssd1 vccd1 vccd1 _19551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16763_ _16761_/X _19312_/Q _16775_/S vssd1 vssd1 vccd1 vccd1 _16764_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13975_ _13975_/A vssd1 vssd1 vccd1 vccd1 _13975_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15713__S _15719_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18502_ _19079_/CLK _18502_/D vssd1 vssd1 vccd1 vccd1 _18502_/Q sky130_fd_sc_hd__dfxtp_2
X_15714_ _15714_/A vssd1 vssd1 vccd1 vccd1 _18870_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12926_ _18286_/Q _12926_/B _12926_/C vssd1 vssd1 vccd1 vccd1 _12933_/D sky130_fd_sc_hd__and3_1
X_19482_ _19682_/CLK _19482_/D vssd1 vssd1 vccd1 vccd1 _19482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16694_ _19291_/Q _16693_/X _16703_/S vssd1 vssd1 vccd1 vccd1 _16695_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18433_ _19695_/CLK _18433_/D vssd1 vssd1 vccd1 vccd1 _18433_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15776__A0 _14918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15645_ _18840_/Q _15564_/X _15647_/S vssd1 vssd1 vccd1 vccd1 _15646_/A sky130_fd_sc_hd__mux2_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12857_ _18266_/Q _12851_/C _12856_/Y vssd1 vssd1 vccd1 vccd1 _18266_/D sky130_fd_sc_hd__o21a_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18364_ _18381_/CLK _18364_/D vssd1 vssd1 vccd1 vccd1 _18364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11808_ _13984_/A _11808_/B vssd1 vssd1 vccd1 vccd1 _11810_/A sky130_fd_sc_hd__xnor2_4
XFILLER_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12788_ _18553_/Q _18552_/Q _18536_/Q _18535_/Q vssd1 vssd1 vccd1 vccd1 _12789_/D
+ sky130_fd_sc_hd__or4_1
X_15576_ _15576_/A vssd1 vssd1 vccd1 vccd1 _18811_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _19531_/Q _16737_/X _17317_/S vssd1 vssd1 vccd1 vccd1 _17316_/A sky130_fd_sc_hd__mux2_1
X_14527_ _11511_/A _12763_/X _14526_/Y _14514_/X vssd1 vssd1 vccd1 vccd1 _18529_/D
+ sky130_fd_sc_hd__o211a_1
X_11739_ _12465_/A _11738_/Y _12173_/A vssd1 vssd1 vccd1 vccd1 _11740_/A sky130_fd_sc_hd__mux2_2
X_18295_ _18298_/CLK _18295_/D vssd1 vssd1 vccd1 vccd1 _18295_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18190__A1 _19850_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17246_ _17246_/A vssd1 vssd1 vccd1 vccd1 _19500_/D sky130_fd_sc_hd__clkbuf_1
X_14458_ _14458_/A vssd1 vssd1 vccd1 vccd1 _18500_/D sky130_fd_sc_hd__clkbuf_1
X_13409_ _18332_/Q _13178_/X _12665_/A _19821_/Q _13408_/X vssd1 vssd1 vccd1 vccd1
+ _13409_/X sky130_fd_sc_hd__a221o_1
XANTENNA__14751__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17177_ _17177_/A vssd1 vssd1 vccd1 vccd1 _19479_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14751__B2 _14711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14389_ _18475_/Q vssd1 vssd1 vccd1 vccd1 _17701_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_152_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19568_/CLK sky130_fd_sc_hd__clkbuf_16
X_16128_ _16838_/A vssd1 vssd1 vccd1 vccd1 _16128_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16059_ _16058_/X _19021_/Q _16065_/S vssd1 vssd1 vccd1 vccd1 _16060_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_167_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19062_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19818_ _19818_/CLK _19818_/D vssd1 vssd1 vccd1 vccd1 _19818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19749_ _19755_/CLK _19749_/D vssd1 vssd1 vccd1 vccd1 _19749_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16719__S _16719_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17205__A0 _18445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09502_ _10591_/A vssd1 vssd1 vccd1 vccd1 _10227_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15623__S _15625_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17404__A _17461_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09433_ _11205_/A _12505_/A vssd1 vssd1 vccd1 vccd1 _11284_/B sky130_fd_sc_hd__or2_1
XFILLER_53_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ _09364_/A vssd1 vssd1 vccd1 vccd1 _09370_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_105_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _18298_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12267__B _19751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09295_ _18577_/Q vssd1 vssd1 vccd1 vccd1 _14570_/A sky130_fd_sc_hd__inv_2
XANTENNA__18181__A1 _19847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10068__A _10068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11100__S0 _10350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17285__S _17291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_108_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15594__A _15662_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput160 _12301_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[24] sky130_fd_sc_hd__buf_2
XFILLER_88_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput171 _11804_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[5] sky130_fd_sc_hd__buf_2
XFILLER_88_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09592__A _09675_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10070_ _10064_/A _10069_/X _09318_/A vssd1 vssd1 vccd1 vccd1 _10070_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15533__S _15536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13760_ _13756_/X _13955_/B _13991_/S vssd1 vssd1 vccd1 vccd1 _13760_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10972_ _19406_/Q _19182_/Q _19699_/Q _19150_/Q _10919_/X _10920_/X vssd1 vssd1 vccd1
+ vccd1 _10973_/B sky130_fd_sc_hd__mux4_1
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12711_ _18630_/Q _12711_/B vssd1 vssd1 vccd1 vccd1 _12711_/X sky130_fd_sc_hd__or2_1
XFILLER_16_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13691_ _13687_/X _13690_/X _13759_/S vssd1 vssd1 vccd1 vccd1 _13691_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12458__A _12458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12642_ _12642_/A vssd1 vssd1 vccd1 vccd1 _13127_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15430_ _15430_/A vssd1 vssd1 vccd1 vccd1 _18758_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15361_ _15361_/A vssd1 vssd1 vccd1 vccd1 _18729_/D sky130_fd_sc_hd__clkbuf_1
X_12573_ _14601_/A vssd1 vssd1 vccd1 vccd1 _17895_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__14981__A1 _12756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14673__A _14673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17100_ _16793_/X _19450_/Q _17108_/S vssd1 vssd1 vccd1 vccd1 _17101_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09767__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14312_ _14312_/A _14312_/B vssd1 vssd1 vccd1 vccd1 _14312_/X sky130_fd_sc_hd__or2_1
X_11524_ _11692_/B vssd1 vssd1 vccd1 vccd1 _12466_/B sky130_fd_sc_hd__buf_2
X_18080_ _18114_/A _18086_/C vssd1 vssd1 vccd1 vccd1 _18080_/Y sky130_fd_sc_hd__nor2_1
X_15292_ _18699_/Q _15171_/X _15300_/S vssd1 vssd1 vccd1 vccd1 _15293_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15488__B _16357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14243_ _14003_/X _14240_/Y _14242_/X vssd1 vssd1 vccd1 vccd1 _14243_/Y sky130_fd_sc_hd__o21ai_1
X_17031_ _17031_/A vssd1 vssd1 vccd1 vccd1 _19419_/D sky130_fd_sc_hd__clkbuf_1
X_11455_ _14426_/A vssd1 vssd1 vccd1 vccd1 _14120_/A sky130_fd_sc_hd__buf_2
XANTENNA__12193__A _17143_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10406_ _19643_/Q _19060_/Q _19097_/Q _18703_/Q _09673_/S _09602_/A vssd1 vssd1 vccd1
+ vccd1 _10406_/X sky130_fd_sc_hd__mux4_1
X_14174_ _13909_/X _14171_/X _14172_/Y _15123_/A vssd1 vssd1 vccd1 vccd1 _14174_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_109_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11386_ _18427_/Q _18426_/Q _11306_/X _11385_/Y vssd1 vssd1 vccd1 vccd1 _11722_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_124_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13125_ _19469_/Q _13203_/A _13205_/A _18383_/Q vssd1 vssd1 vccd1 vccd1 _13125_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15708__S _15708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_84_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19496_/CLK sky130_fd_sc_hd__clkbuf_16
X_10337_ _11185_/A _10337_/B vssd1 vssd1 vccd1 vccd1 _10337_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18982_ _18982_/CLK _18982_/D vssd1 vssd1 vccd1 vccd1 _18982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _17934_/B _17934_/C _19763_/Q vssd1 vssd1 vccd1 vccd1 _17935_/B sky130_fd_sc_hd__a21oi_1
X_13056_ _17935_/A _13056_/B _13056_/C vssd1 vssd1 vccd1 vccd1 _18329_/D sky130_fd_sc_hd__nor3_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10268_ _09995_/A _10267_/X _09214_/A vssd1 vssd1 vccd1 vccd1 _10268_/X sky130_fd_sc_hd__o21a_1
XFILLER_140_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09912__A1 _09149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12007_ _14089_/B _11972_/B _12106_/A vssd1 vssd1 vccd1 vccd1 _12008_/B sky130_fd_sc_hd__a21o_1
X_17864_ _11803_/A _11803_/B _14638_/A vssd1 vssd1 vccd1 vccd1 _19733_/D sky130_fd_sc_hd__a21o_1
XFILLER_39_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10199_ _10212_/A _10199_/B vssd1 vssd1 vccd1 vccd1 _10199_/X sky130_fd_sc_hd__or2_1
XFILLER_78_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_99_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19690_/CLK sky130_fd_sc_hd__clkbuf_16
X_19603_ _19702_/CLK _19603_/D vssd1 vssd1 vccd1 vccd1 _19603_/Q sky130_fd_sc_hd__dfxtp_1
X_16815_ _16815_/A vssd1 vssd1 vccd1 vccd1 _19328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17795_ _17795_/A vssd1 vssd1 vccd1 vccd1 _19700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16539__S _16547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19534_ _19534_/CLK _19534_/D vssd1 vssd1 vccd1 vccd1 _19534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16746_ _16845_/S vssd1 vssd1 vccd1 vccd1 _16759_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_59_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13958_ _13838_/A _13954_/X _13957_/Y _14036_/S vssd1 vssd1 vccd1 vccd1 _13958_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_46_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10286__A1 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12909_ _18281_/Q _12907_/B _12908_/Y vssd1 vssd1 vccd1 vccd1 _18281_/D sky130_fd_sc_hd__o21a_1
X_19465_ _19595_/CLK _19465_/D vssd1 vssd1 vccd1 vccd1 _19465_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_22_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19714_/CLK sky130_fd_sc_hd__clkbuf_16
X_16677_ _16677_/A vssd1 vssd1 vccd1 vccd1 _16677_/X sky130_fd_sc_hd__buf_2
XFILLER_61_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12368__A _13388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13889_ _13774_/Y _13887_/Y _13888_/X _13913_/S vssd1 vssd1 vccd1 vccd1 _13889_/X
+ sky130_fd_sc_hd__a22o_1
X_18416_ _19481_/CLK _18416_/D vssd1 vssd1 vccd1 vccd1 _18416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15628_ _18832_/Q _15538_/X _15636_/S vssd1 vssd1 vccd1 vccd1 _15629_/A sky130_fd_sc_hd__mux2_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19396_ _19590_/CLK _19396_/D vssd1 vssd1 vccd1 vccd1 _19396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18347_ _19759_/CLK _18347_/D vssd1 vssd1 vccd1 vccd1 _18347_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09523__S0 _11110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14972__A1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15559_ _18806_/Q _15558_/X _15568_/S vssd1 vssd1 vccd1 vccd1 _15560_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_37_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19626_/CLK sky130_fd_sc_hd__clkbuf_16
X_09080_ _09125_/A _18567_/Q vssd1 vssd1 vccd1 vccd1 _09107_/A sky130_fd_sc_hd__or2_1
X_18278_ _18401_/CLK _18278_/D vssd1 vssd1 vccd1 vccd1 _18278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput40 io_ibus_inst[15] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_2
X_17229_ _18452_/Q _13376_/X _17235_/S vssd1 vssd1 vccd1 vccd1 _17229_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput51 io_ibus_inst[25] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_2
XANTENNA__10616__A _10906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput62 io_ibus_inst[6] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09982_ _10256_/S vssd1 vssd1 vccd1 vccd1 _10200_/S sky130_fd_sc_hd__buf_4
XFILLER_104_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09416_ _19628_/Q _19466_/Q _18912_/Q _18682_/Q _09367_/S _09364_/A vssd1 vssd1 vccd1
+ vccd1 _09417_/B sky130_fd_sc_hd__mux4_1
XFILLER_80_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_34_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09347_ _09955_/A vssd1 vssd1 vccd1 vccd1 _09928_/A sky130_fd_sc_hd__buf_4
XANTENNA__18154__A1 _19838_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09587__A _09587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09278_ _09278_/A vssd1 vssd1 vccd1 vccd1 _09278_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_166_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13518__A2 _12731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_3_0_clock_A clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11240_ _11262_/A _11262_/B vssd1 vssd1 vccd1 vccd1 _11263_/A sky130_fd_sc_hd__and2_1
XFILLER_134_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17665__A0 _19670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11171_ _11171_/A _11171_/B vssd1 vssd1 vccd1 vccd1 _11171_/X sky130_fd_sc_hd__or2_1
XANTENNA__12741__A _13235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16213__A _17783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10122_ _10020_/A _10121_/X _09988_/X vssd1 vssd1 vccd1 vccd1 _10122_/X sky130_fd_sc_hd__o21a_1
XFILLER_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18209__A2 _18214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12460__B _12466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10053_ _18869_/Q _19327_/Q _10055_/S vssd1 vssd1 vccd1 vccd1 _10054_/B sky130_fd_sc_hd__mux2_1
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14930_ _14929_/X _18604_/Q _14941_/S vssd1 vssd1 vccd1 vccd1 _14931_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15979__A0 _14792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A io_dbus_rdata[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861_ _14861_/A _18471_/Q _14861_/C vssd1 vssd1 vccd1 vccd1 _14871_/B sky130_fd_sc_hd__and3_1
XFILLER_29_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16600_ _16600_/A vssd1 vssd1 vccd1 vccd1 _19255_/D sky130_fd_sc_hd__clkbuf_1
X_13812_ _13811_/Y _13703_/A _13880_/S vssd1 vssd1 vccd1 vccd1 _13812_/X sky130_fd_sc_hd__mux2_1
X_17580_ _17580_/A vssd1 vssd1 vccd1 vccd1 _19648_/D sky130_fd_sc_hd__clkbuf_1
X_14792_ _16768_/A vssd1 vssd1 vccd1 vccd1 _14792_/X sky130_fd_sc_hd__buf_2
XANTENNA__12257__A2 _14227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16531_ _16531_/A vssd1 vssd1 vccd1 vccd1 _19222_/D sky130_fd_sc_hd__clkbuf_1
X_13743_ _13741_/X _13742_/X _13743_/S vssd1 vssd1 vccd1 vccd1 _13743_/X sky130_fd_sc_hd__mux2_1
X_10955_ _18820_/Q _19374_/Q _19536_/Q _18788_/Q _10909_/X _10910_/X vssd1 vssd1 vccd1
+ vccd1 _10956_/B sky130_fd_sc_hd__mux4_1
XFILLER_73_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12188__A _19748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19250_ _19634_/CLK _19250_/D vssd1 vssd1 vccd1 vccd1 _19250_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13206__A1 _19665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16462_ _16077_/X _19192_/Q _16464_/S vssd1 vssd1 vccd1 vccd1 _16463_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10200__S _10200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13674_ _13776_/S vssd1 vssd1 vccd1 vccd1 _13877_/S sky130_fd_sc_hd__clkbuf_2
X_10886_ _18588_/Q _19277_/Q _10886_/S vssd1 vssd1 vccd1 vccd1 _10887_/B sky130_fd_sc_hd__mux2_1
XFILLER_71_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18201_ _18223_/A _18201_/B vssd1 vssd1 vccd1 vccd1 _18201_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15413_ _15413_/A _15960_/C vssd1 vssd1 vccd1 vccd1 _16992_/A sky130_fd_sc_hd__or2_4
XANTENNA__09505__S0 _10277_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12625_ _18344_/Q _12643_/A _12669_/A _19488_/Q vssd1 vssd1 vccd1 vccd1 _12625_/X
+ sky130_fd_sc_hd__a22o_1
X_19181_ _19633_/CLK _19181_/D vssd1 vssd1 vccd1 vccd1 _19181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16393_ _16415_/A vssd1 vssd1 vccd1 vccd1 _16402_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__16094__S _16097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18132_ _18165_/A _18132_/B _18132_/C vssd1 vssd1 vccd1 vccd1 _19830_/D sky130_fd_sc_hd__nor3_1
XANTENNA__09497__A _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12556_ _12600_/A vssd1 vssd1 vccd1 vccd1 _12556_/X sky130_fd_sc_hd__buf_2
X_15344_ _15344_/A vssd1 vssd1 vccd1 vccd1 _18721_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11507_ _15079_/A _13527_/B _13529_/A vssd1 vssd1 vccd1 vccd1 _11508_/C sky130_fd_sc_hd__and3_1
XFILLER_156_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18063_ _18071_/A _18067_/C vssd1 vssd1 vccd1 vccd1 _18063_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15275_ _15275_/A vssd1 vssd1 vccd1 vccd1 _18691_/D sky130_fd_sc_hd__clkbuf_1
X_12487_ _12487_/A _12497_/B vssd1 vssd1 vccd1 vccd1 _12487_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17014_ _19412_/Q _16670_/X _17014_/S vssd1 vssd1 vccd1 vccd1 _17015_/A sky130_fd_sc_hd__mux2_1
X_11438_ _12557_/A _11438_/B vssd1 vssd1 vccd1 vccd1 _13108_/B sky130_fd_sc_hd__nor2_4
X_14226_ _14088_/X _14223_/Y _14225_/X vssd1 vssd1 vccd1 vccd1 _14226_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_160_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14157_ _13788_/A _14154_/X _14156_/Y _13894_/A vssd1 vssd1 vccd1 vccd1 _14157_/X
+ sky130_fd_sc_hd__a31o_1
X_11369_ _11692_/A _11592_/A _11593_/A _11368_/X vssd1 vssd1 vccd1 vccd1 _11369_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_140_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09686__A1_N _18453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13108_ _13108_/A _13108_/B vssd1 vssd1 vccd1 vccd1 _13442_/D sky130_fd_sc_hd__nor2_1
XANTENNA__15131__A1 _18649_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18965_ _19295_/CLK _18965_/D vssd1 vssd1 vccd1 vccd1 _18965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ _14088_/A vssd1 vssd1 vccd1 vccd1 _14088_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15131__B2 _11202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13039_ _18325_/Q vssd1 vssd1 vccd1 vccd1 _13045_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17916_ _19803_/Q _19802_/Q _19804_/Q _18046_/A vssd1 vssd1 vccd1 vccd1 _18054_/A
+ sky130_fd_sc_hd__and4_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18896_ _19551_/CLK _18896_/D vssd1 vssd1 vccd1 vccd1 _18896_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09960__A _09969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17847_ _15229_/X _19724_/Q _17849_/S vssd1 vssd1 vccd1 vccd1 _17848_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14578__A _14578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15173__S _15185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13445__A1 _13136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17778_ _17778_/A vssd1 vssd1 vccd1 vccd1 _19693_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19517_ _19612_/CLK _19517_/D vssd1 vssd1 vccd1 vccd1 _19517_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11456__A0 _14737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09744__S0 _09721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16729_ _19302_/Q _16728_/X _16735_/S vssd1 vssd1 vccd1 vccd1 _16730_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12098__A _19675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16793__A _16793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19448_ _19610_/CLK _19448_/D vssd1 vssd1 vccd1 vccd1 _19448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09201_ _10313_/A vssd1 vssd1 vccd1 vccd1 _10212_/A sky130_fd_sc_hd__buf_2
XFILLER_50_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19379_ _19539_/CLK _19379_/D vssd1 vssd1 vccd1 vccd1 _19379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10106__S1 _10103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09132_ _10373_/A vssd1 vssd1 vccd1 vccd1 _09133_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_136_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09200__A _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16732__S _16735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17647__A0 _19667_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12561__A _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09965_ _09969_/A _09965_/B vssd1 vssd1 vccd1 vccd1 _09965_/X sky130_fd_sc_hd__or2_1
XANTENNA__15122__B2 _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09896_ _18451_/Q _09309_/X _09430_/X _09895_/X vssd1 vssd1 vccd1 vccd1 _12499_/A
+ sky130_fd_sc_hd__o2bb2a_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16179__S _16183_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_10_0_clock_A clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16907__S _16913_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15811__S _15819_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10740_ _10740_/A vssd1 vssd1 vccd1 vccd1 _10740_/X sky130_fd_sc_hd__buf_2
XANTENNA__15189__A1 _15187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ _10605_/S _10666_/Y _10669_/Y _10670_/X vssd1 vssd1 vccd1 vccd1 _10671_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_41_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ _19757_/Q _12410_/B vssd1 vssd1 vccd1 vccd1 _12411_/C sky130_fd_sc_hd__or2_1
XFILLER_139_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13390_ _13390_/A _18647_/Q vssd1 vssd1 vccd1 vccd1 _13390_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09812__B1 _09415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12341_ _18376_/Q _12341_/B vssd1 vssd1 vccd1 vccd1 _12393_/C sky130_fd_sc_hd__and2_1
XANTENNA__14663__A1_N input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15060_ _18456_/Q _15060_/B vssd1 vssd1 vccd1 vccd1 _15060_/X sky130_fd_sc_hd__or2_1
X_12272_ _18373_/Q _18372_/Q _12272_/C vssd1 vssd1 vccd1 vccd1 _12320_/C sky130_fd_sc_hd__and3_1
XFILLER_107_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14011_ _14000_/X _14002_/X _14010_/Y _13594_/A vssd1 vssd1 vccd1 vccd1 _14011_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11223_ _09756_/B _11221_/X _11222_/X vssd1 vssd1 vccd1 vccd1 _11223_/X sky130_fd_sc_hd__a21o_1
XFILLER_134_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11154_ _19271_/Q _19042_/Q _18973_/Q _19367_/Q _11153_/X _10306_/X vssd1 vssd1 vccd1
+ vccd1 _11155_/B sky130_fd_sc_hd__mux4_1
XFILLER_108_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15113__B2 _10299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7_0_clock_A clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10105_ _10120_/A _10105_/B vssd1 vssd1 vccd1 vccd1 _10105_/X sky130_fd_sc_hd__or2_1
X_18750_ _19725_/CLK _18750_/D vssd1 vssd1 vccd1 vccd1 _18750_/Q sky130_fd_sc_hd__dfxtp_1
X_15962_ _16018_/A vssd1 vssd1 vccd1 vccd1 _16031_/S sky130_fd_sc_hd__buf_8
X_11085_ _19256_/Q _19027_/Q _18958_/Q _19352_/Q _09447_/A _09635_/A vssd1 vssd1 vccd1
+ vccd1 _11086_/B sky130_fd_sc_hd__mux4_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09780__A _10094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17701_ _17701_/A _17701_/B _17701_/C vssd1 vssd1 vccd1 vccd1 _17710_/B sky130_fd_sc_hd__or3_1
X_10036_ _18774_/Q _19003_/Q _18934_/Q _19232_/Q _09866_/A _10029_/X vssd1 vssd1 vccd1
+ vccd1 _10037_/B sky130_fd_sc_hd__mux4_1
XFILLER_76_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14913_ _17701_/A _14912_/B _14945_/B vssd1 vssd1 vccd1 vccd1 _14913_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_102_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18681_ _19726_/CLK _18681_/D vssd1 vssd1 vccd1 vccd1 _18681_/Q sky130_fd_sc_hd__dfxtp_1
X_15893_ _15950_/S vssd1 vssd1 vccd1 vccd1 _15902_/S sky130_fd_sc_hd__buf_4
XFILLER_36_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11815__A _11849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17632_ _17632_/A _18464_/Q _17632_/C vssd1 vssd1 vccd1 vccd1 _17640_/B sky130_fd_sc_hd__or3_1
XFILLER_75_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14844_ _14838_/X _14839_/X _14843_/Y vssd1 vssd1 vccd1 vccd1 _14845_/B sky130_fd_sc_hd__a21oi_4
XFILLER_90_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17563_ _17563_/A vssd1 vssd1 vccd1 vccd1 _19640_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14775_ _14775_/A vssd1 vssd1 vccd1 vccd1 _18591_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16817__S _16823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11987_ _11978_/X _11985_/Y _12294_/S vssd1 vssd1 vccd1 vccd1 _11987_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19302_ _19624_/CLK _19302_/D vssd1 vssd1 vccd1 vccd1 _19302_/Q sky130_fd_sc_hd__dfxtp_1
X_16514_ _19215_/Q _15503_/X _16514_/S vssd1 vssd1 vccd1 vccd1 _16515_/A sky130_fd_sc_hd__mux2_1
X_13726_ _13950_/A vssd1 vssd1 vccd1 vccd1 _13726_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10938_ _19406_/Q _19182_/Q _19699_/Q _19150_/Q _10706_/S _09352_/A vssd1 vssd1 vccd1
+ vccd1 _10938_/X sky130_fd_sc_hd__mux4_1
X_17494_ _19610_/Q _16683_/X _17496_/S vssd1 vssd1 vccd1 vccd1 _17495_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19233_ _19555_/CLK _19233_/D vssd1 vssd1 vccd1 vccd1 _19233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16445_ _16051_/X _19184_/Q _16453_/S vssd1 vssd1 vccd1 vccd1 _16446_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14927__A1 _11542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13657_ _14265_/B _13984_/B _13657_/S vssd1 vssd1 vccd1 vccd1 _13657_/X sky130_fd_sc_hd__mux2_1
X_10869_ _10827_/X _10866_/Y _10868_/Y _09244_/A vssd1 vssd1 vccd1 vccd1 _10869_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_32_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12938__B1 _18290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12608_ _18345_/Q _12643_/A _12539_/A _19677_/Q vssd1 vssd1 vccd1 vccd1 _12608_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19164_ _19713_/CLK _19164_/D vssd1 vssd1 vccd1 vccd1 _19164_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _19154_/Q _15513_/X _16380_/S vssd1 vssd1 vccd1 vccd1 _16377_/A sky130_fd_sc_hd__mux2_1
X_13588_ _13720_/B vssd1 vssd1 vccd1 vccd1 _13729_/B sky130_fd_sc_hd__clkbuf_2
X_18115_ _19825_/Q _18111_/C _18114_/Y vssd1 vssd1 vccd1 vccd1 _19825_/D sky130_fd_sc_hd__o21a_1
XFILLER_9_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15327_ _18715_/Q _15223_/X _15333_/S vssd1 vssd1 vccd1 vccd1 _15328_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15957__A _15957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12539_ _12539_/A vssd1 vssd1 vccd1 vccd1 _12624_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16552__S _16558_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19095_ _19579_/CLK _19095_/D vssd1 vssd1 vccd1 vccd1 _19095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18046_ _18046_/A vssd1 vssd1 vccd1 vccd1 _18051_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15258_ _15262_/A vssd1 vssd1 vccd1 vccd1 _15258_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14209_ _18446_/Q _14208_/X _14209_/S vssd1 vssd1 vccd1 vccd1 _14210_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12381__A _12381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15189_ _18666_/Q _15187_/X _15201_/S vssd1 vssd1 vccd1 vccd1 _15190_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13196__B _13196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17383__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09750_ _09743_/Y _09745_/Y _09747_/Y _09749_/Y _09403_/A vssd1 vssd1 vccd1 vccd1
+ _09750_/X sky130_fd_sc_hd__o221a_2
X_18948_ _19631_/CLK _18948_/D vssd1 vssd1 vccd1 vccd1 _18948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11126__C1 _10494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10024__S0 _10076_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09690__A _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09681_ _09681_/A vssd1 vssd1 vccd1 vccd1 _09681_/X sky130_fd_sc_hd__buf_2
XFILLER_95_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18879_ _19337_/CLK _18879_/D vssd1 vssd1 vccd1 vccd1 _18879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17801__A0 _15162_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10575__S1 _10368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15040__A0 _18454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12556__A _12600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12929__B1 _18287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09115_ _18566_/Q vssd1 vssd1 vccd1 vccd1 _11343_/B sky130_fd_sc_hd__inv_2
XFILLER_129_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16462__S _16464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15343__A1 _15133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12291__A _19752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15806__S _15806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09948_ _09944_/A _09945_/X _09947_/X _09320_/A vssd1 vssd1 vccd1 vccd1 _09948_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_77_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10015__S0 _10076_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09879_ _09879_/A vssd1 vssd1 vccd1 vccd1 _09944_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _19737_/Q _11705_/X _11905_/X _11909_/X vssd1 vssd1 vccd1 vccd1 _17872_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_85_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10340__A0 _19612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12890_ _12895_/C _12893_/C _12869_/X vssd1 vssd1 vccd1 vccd1 _12890_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11354__B _11514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _10691_/X _18497_/Q _11948_/A vssd1 vssd1 vccd1 vccd1 _13658_/A sky130_fd_sc_hd__mux2_8
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14946__A _14958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10318__S1 _10306_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _11756_/X _11771_/Y _19732_/Q _11788_/B vssd1 vssd1 vccd1 vccd1 _17862_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14560_ _14585_/A vssd1 vssd1 vccd1 vccd1 _14560_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _13511_/A vssd1 vssd1 vccd1 vccd1 _18413_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10643__A1 _09409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10723_ _10797_/A vssd1 vssd1 vccd1 vccd1 _10803_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14491_ _14491_/A vssd1 vssd1 vccd1 vccd1 _18515_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12466__A _12466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16230_ _16230_/A vssd1 vssd1 vccd1 vccd1 _19089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13442_ _12541_/B _12791_/B _13442_/C _13442_/D vssd1 vssd1 vccd1 vccd1 _13499_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_110_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10654_ _19411_/Q _19187_/Q _19704_/Q _19155_/Q _10836_/A _09353_/A vssd1 vssd1 vccd1
+ vccd1 _10654_/X sky130_fd_sc_hd__mux4_1
XFILLER_167_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17468__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12396__B2 _12503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13373_ _19850_/Q _12736_/X _13371_/X _13372_/X vssd1 vssd1 vccd1 vccd1 _13373_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17859__B1 _14638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16161_ _16064_/X _19055_/Q _16161_/S vssd1 vssd1 vccd1 vccd1 _16162_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10585_ _19412_/Q _19188_/Q _19705_/Q _19156_/Q _10511_/S _09662_/A vssd1 vssd1 vccd1
+ vccd1 _10585_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15112_ _18634_/Q _15109_/X _15111_/X _11135_/A vssd1 vssd1 vccd1 vccd1 _18634_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_155_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12324_ _14578_/A _12344_/A _12345_/A _12500_/A vssd1 vssd1 vccd1 vccd1 _12325_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_16092_ _16092_/A vssd1 vssd1 vccd1 vccd1 _19031_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15043_ _16731_/A vssd1 vssd1 vccd1 vccd1 _16835_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12255_ _12495_/C _12345_/A _12254_/X vssd1 vssd1 vccd1 vccd1 _12256_/A sky130_fd_sc_hd__o21ai_1
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_3_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11206_ _11203_/A _11204_/Y _11205_/Y _11284_/B vssd1 vssd1 vccd1 vccd1 _11207_/A
+ sky130_fd_sc_hd__o211ai_1
X_19851_ _19851_/CLK _19851_/D vssd1 vssd1 vccd1 vccd1 _19851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12186_ _12186_/A vssd1 vssd1 vccd1 vccd1 _12186_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_156_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18802_ _19713_/CLK _18802_/D vssd1 vssd1 vccd1 vccd1 _18802_/Q sky130_fd_sc_hd__dfxtp_1
X_11137_ _11137_/A _12486_/A vssd1 vssd1 vccd1 vccd1 _11137_/X sky130_fd_sc_hd__and2_1
XFILLER_95_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19782_ _19861_/CLK _19782_/D vssd1 vssd1 vccd1 vccd1 _19782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16994_ _17062_/S vssd1 vssd1 vccd1 vccd1 _17003_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_62_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18733_ _19708_/CLK _18733_/D vssd1 vssd1 vccd1 vccd1 _18733_/Q sky130_fd_sc_hd__dfxtp_1
X_15945_ _15945_/A vssd1 vssd1 vccd1 vccd1 _18973_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11068_ _09926_/A _11058_/X _11067_/X _09305_/A _11046_/A vssd1 vssd1 vccd1 vccd1
+ _12458_/A sky130_fd_sc_hd__a32o_4
XFILLER_37_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10019_ _19650_/Q _19067_/Q _19104_/Q _18710_/Q _09782_/A _09979_/X vssd1 vssd1 vccd1
+ vccd1 _10020_/B sky130_fd_sc_hd__mux4_1
XFILLER_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18664_ _19610_/CLK _18664_/D vssd1 vssd1 vccd1 vccd1 _18664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15876_ _15066_/X _18943_/Q _15878_/S vssd1 vssd1 vccd1 vccd1 _15877_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17615_ _19661_/Q _17610_/X _17625_/S vssd1 vssd1 vccd1 vccd1 _17616_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14827_ _18467_/Q _18468_/Q _14827_/C vssd1 vssd1 vccd1 vccd1 _14840_/B sky130_fd_sc_hd__and3_1
X_18595_ _19444_/CLK _18595_/D vssd1 vssd1 vccd1 vccd1 _18595_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16547__S _16547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14856__A _16784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15451__S _15459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17546_ _19633_/Q _16758_/A _17546_/S vssd1 vssd1 vccd1 vccd1 _17547_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14758_ _14756_/X _14757_/X _14923_/S vssd1 vssd1 vccd1 vccd1 _14758_/X sky130_fd_sc_hd__mux2_2
XFILLER_149_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13709_ _14276_/A vssd1 vssd1 vccd1 vccd1 _14312_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17477_ _19602_/Q _16657_/X _17485_/S vssd1 vssd1 vccd1 vccd1 _17478_/A sky130_fd_sc_hd__mux2_1
X_14689_ _14689_/A vssd1 vssd1 vccd1 vccd1 _18582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19216_ _19569_/CLK _19216_/D vssd1 vssd1 vccd1 vccd1 _19216_/Q sky130_fd_sc_hd__dfxtp_1
X_16428_ _19178_/Q _15589_/X _16428_/S vssd1 vssd1 vccd1 vccd1 _16429_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19147_ _19436_/CLK _19147_/D vssd1 vssd1 vccd1 vccd1 _19147_/Q sky130_fd_sc_hd__dfxtp_1
X_16359_ _16415_/A vssd1 vssd1 vccd1 vccd1 _16428_/S sky130_fd_sc_hd__buf_8
XFILLER_146_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19078_ _19078_/CLK _19078_/D vssd1 vssd1 vccd1 vccd1 _19078_/Q sky130_fd_sc_hd__dfxtp_1
X_18029_ _18031_/B _18031_/C _17993_/X vssd1 vssd1 vccd1 vccd1 _18029_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_161_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11439__B _18417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15089__A0 _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09802_ _10033_/S vssd1 vssd1 vccd1 vccd1 _09803_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10796__S1 _10713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09733_ _11185_/A vssd1 vssd1 vccd1 vccd1 _10127_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17841__S _17849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09664_ _10390_/A vssd1 vssd1 vccd1 vccd1 _10280_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17250__A1 _16639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09595_ _09595_/A _09595_/B vssd1 vssd1 vccd1 vccd1 _09595_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12286__A _12286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10720__S1 _09481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16192__S _16194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09595__A _09595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10370_ _18767_/Q _18996_/Q _18927_/Q _19225_/Q _09631_/A _10368_/A vssd1 vssd1 vccd1
+ vccd1 _10371_/B sky130_fd_sc_hd__mux4_1
XFILLER_163_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12040_ _12040_/A _12040_/B vssd1 vssd1 vccd1 vccd1 _12041_/A sky130_fd_sc_hd__xnor2_4
XFILLER_85_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10253__B _12486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15536__S _15536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13991_ _13876_/X _13879_/X _13991_/S vssd1 vssd1 vccd1 vccd1 _13992_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11105__A2 _11095_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12302__B2 _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15730_ _18878_/Q _15583_/X _15730_/S vssd1 vssd1 vccd1 vccd1 _15731_/A sky130_fd_sc_hd__mux2_1
X_12942_ _18291_/Q _12946_/C vssd1 vssd1 vccd1 vccd1 _12945_/B sky130_fd_sc_hd__and2_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17241__A1 _13423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _15661_/A vssd1 vssd1 vccd1 vccd1 _18847_/D sky130_fd_sc_hd__clkbuf_1
X_12873_ _18271_/Q _12873_/B _12873_/C vssd1 vssd1 vccd1 vccd1 _12874_/C sky130_fd_sc_hd__and3_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16367__S _16369_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _16755_/X _19568_/Q _17402_/S vssd1 vssd1 vccd1 vccd1 _17401_/A sky130_fd_sc_hd__mux2_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _14612_/A _14612_/B vssd1 vssd1 vccd1 vccd1 _18558_/D sky130_fd_sc_hd__nand2_1
X_11824_ _11798_/Y _11822_/X _11823_/Y vssd1 vssd1 vccd1 vccd1 _11826_/B sky130_fd_sc_hd__a21o_1
X_18380_ _18381_/CLK _18380_/D vssd1 vssd1 vccd1 vccd1 _18380_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _16992_/A _15592_/B vssd1 vssd1 vccd1 vccd1 _15649_/A sky130_fd_sc_hd__nor2_2
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17331_/A vssd1 vssd1 vccd1 vccd1 _19537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14543_ _14543_/A _14551_/B vssd1 vssd1 vccd1 vccd1 _14543_/Y sky130_fd_sc_hd__nand2_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12196__A _17628_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11755_ _19663_/Q _12412_/B _17221_/A vssd1 vssd1 vccd1 vccd1 _11755_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15004__B1 _14737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_82_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10706_ _18593_/Q _19282_/Q _10706_/S vssd1 vssd1 vccd1 vccd1 _10706_/X sky130_fd_sc_hd__mux2_1
X_17262_ _17262_/A vssd1 vssd1 vccd1 vccd1 _19506_/D sky130_fd_sc_hd__clkbuf_1
X_14474_ _18508_/Q _19746_/Q _14476_/S vssd1 vssd1 vccd1 vccd1 _14475_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11686_ _11686_/A _11686_/B _13587_/B _11686_/D vssd1 vssd1 vccd1 vccd1 _11776_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_174_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19001_ _19326_/CLK _19001_/D vssd1 vssd1 vccd1 vccd1 _19001_/Q sky130_fd_sc_hd__dfxtp_1
X_16213_ _17783_/A _16213_/B vssd1 vssd1 vccd1 vccd1 _16270_/A sky130_fd_sc_hd__nand2_2
X_13425_ _13311_/A _13423_/X _13424_/X _13401_/X vssd1 vssd1 vccd1 vccd1 _18380_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17193_ _19484_/Q _17191_/X _17206_/S vssd1 vssd1 vccd1 vccd1 _17194_/A sky130_fd_sc_hd__mux2_1
X_10637_ _18825_/Q _19379_/Q _19541_/Q _18793_/Q _10631_/X _10634_/X vssd1 vssd1 vccd1
+ vccd1 _10638_/B sky130_fd_sc_hd__mux4_2
XFILLER_127_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16144_ _16039_/X _19047_/Q _16150_/S vssd1 vssd1 vccd1 vccd1 _16145_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15307__A1 _15194_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13356_ _18292_/Q _12638_/X _13127_/X _18375_/Q vssd1 vssd1 vccd1 vccd1 _13356_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10568_ _10568_/A _10568_/B _10568_/C vssd1 vssd1 vccd1 vccd1 _10568_/X sky130_fd_sc_hd__or3_2
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12307_ _12307_/A vssd1 vssd1 vccd1 vccd1 _14265_/B sky130_fd_sc_hd__buf_2
X_16075_ _16074_/X _19026_/Q _16081_/S vssd1 vssd1 vccd1 vccd1 _16076_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13287_ _19673_/Q _12668_/X _12768_/X _18397_/Q vssd1 vssd1 vccd1 vccd1 _13288_/B
+ sky130_fd_sc_hd__a22o_1
X_10499_ _18828_/Q _19382_/Q _19544_/Q _18796_/Q _10242_/S _10239_/A vssd1 vssd1 vccd1
+ vccd1 _10499_/X sky130_fd_sc_hd__mux4_2
XANTENNA__16830__S _16839_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15026_ _15027_/A _15037_/C vssd1 vssd1 vccd1 vccd1 _15026_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14530__A2 _12763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12238_ _12185_/A _12185_/B _12235_/Y _12237_/Y vssd1 vssd1 vccd1 vccd1 _12240_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_69_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10001__C1 _09249_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15446__S _15448_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19834_ _19851_/CLK _19834_/D vssd1 vssd1 vccd1 vccd1 _19834_/Q sky130_fd_sc_hd__dfxtp_2
X_12169_ _18369_/Q _13316_/A _12169_/C vssd1 vssd1 vccd1 vccd1 _12222_/C sky130_fd_sc_hd__and3_1
XFILLER_122_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19765_ _19858_/CLK _19765_/D vssd1 vssd1 vccd1 vccd1 _19765_/Q sky130_fd_sc_hd__dfxtp_1
X_16977_ _16977_/A vssd1 vssd1 vccd1 vccd1 _16986_/S sky130_fd_sc_hd__buf_4
XFILLER_7_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 io_dbus_rdata[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_2
X_15928_ _15928_/A vssd1 vssd1 vccd1 vccd1 _18965_/D sky130_fd_sc_hd__clkbuf_1
X_18716_ _19592_/CLK _18716_/D vssd1 vssd1 vccd1 vccd1 _18716_/Q sky130_fd_sc_hd__dfxtp_1
X_19696_ _19696_/CLK _19696_/D vssd1 vssd1 vccd1 vccd1 _19696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17232__A1 _13387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18647_ _19727_/CLK _18647_/D vssd1 vssd1 vccd1 vccd1 _18647_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10855__A1 _09409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15859_ _14975_/X _18935_/Q _15863_/S vssd1 vssd1 vccd1 vccd1 _15860_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16277__S _16279_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09380_ _10226_/A vssd1 vssd1 vccd1 vccd1 _09661_/A sky130_fd_sc_hd__buf_2
XFILLER_91_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18578_ _18578_/CLK _18578_/D vssd1 vssd1 vccd1 vccd1 _18578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10607__A1 _09538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17529_ _19626_/Q _16734_/X _17529_/S vssd1 vssd1 vccd1 vccd1 _17530_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10702__S1 _09512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15210__A _16712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17836__S _17838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12780__A1 _12779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13665__A _13665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15356__S _15362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09933__C1 _09892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14809__A0 _14808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15880__A _16847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11185__A _11185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17571__S _17579_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ _19623_/Q _19461_/Q _18907_/Q _18677_/Q _09793_/A _09704_/A vssd1 vssd1 vccd1
+ vccd1 _09717_/B sky130_fd_sc_hd__mux4_1
XFILLER_56_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09647_ _09562_/X _09638_/X _09640_/X _09133_/A _09646_/X vssd1 vssd1 vccd1 vccd1
+ _09647_/X sky130_fd_sc_hd__a311o_4
XFILLER_16_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_104_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09578_ _10182_/A _09578_/B vssd1 vssd1 vccd1 vccd1 _09578_/Y sky130_fd_sc_hd__nor2_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16915__S _16917_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11540_ _09624_/A _11460_/X _11539_/X vssd1 vssd1 vccd1 vccd1 _19078_/D sky130_fd_sc_hd__o21a_1
XFILLER_50_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11471_ _11471_/A vssd1 vssd1 vccd1 vccd1 _12495_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13210_ _19475_/Q _13203_/X _13204_/X _13206_/X _13209_/X vssd1 vssd1 vccd1 vccd1
+ _13211_/B sky130_fd_sc_hd__a2111o_2
XANTENNA__12220__A0 _12214_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10422_ _10422_/A vssd1 vssd1 vccd1 vccd1 _10559_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11023__B2 _11022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14190_ _13937_/X _14192_/B _13979_/X _14189_/X vssd1 vssd1 vccd1 vccd1 _14190_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12463__B _12466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13141_ _19470_/Q _13235_/A _13154_/B _18384_/Q vssd1 vssd1 vccd1 vccd1 _13141_/X
+ sky130_fd_sc_hd__a22o_1
X_10353_ _10353_/A vssd1 vssd1 vccd1 vccd1 _10558_/S sky130_fd_sc_hd__buf_2
XFILLER_3_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13278__C _14859_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13072_ _18333_/Q _13068_/C _13071_/Y vssd1 vssd1 vccd1 vccd1 _18333_/D sky130_fd_sc_hd__o21a_1
XFILLER_124_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10209__S0 _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input56_A io_ibus_inst[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14512__A2 _12692_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ _10226_/A _10283_/X _09315_/A vssd1 vssd1 vccd1 vccd1 _10284_/X sky130_fd_sc_hd__o21a_1
XFILLER_151_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16900_ _19362_/Q _16715_/X _16902_/S vssd1 vssd1 vccd1 vccd1 _16901_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12023_ _14589_/A _12023_/B vssd1 vssd1 vccd1 vccd1 _12323_/A sky130_fd_sc_hd__nand2_2
XANTENNA_clkbuf_leaf_29_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17880_ _17882_/A _17880_/B vssd1 vssd1 vccd1 vccd1 _17881_/A sky130_fd_sc_hd__or2_1
Xclkbuf_opt_2_0_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_120_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16831_ _16831_/A vssd1 vssd1 vccd1 vccd1 _19333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17481__S _17485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19550_ _19550_/CLK _19550_/D vssd1 vssd1 vccd1 vccd1 _19550_/Q sky130_fd_sc_hd__dfxtp_1
X_16762_ _16845_/S vssd1 vssd1 vccd1 vccd1 _16775_/S sky130_fd_sc_hd__buf_2
X_13974_ _13974_/A vssd1 vssd1 vccd1 vccd1 _13975_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18501_ _18506_/CLK _18501_/D vssd1 vssd1 vccd1 vccd1 _18501_/Q sky130_fd_sc_hd__dfxtp_1
X_15713_ _18870_/Q _15558_/X _15719_/S vssd1 vssd1 vccd1 vccd1 _15714_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10837__A1 _10631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12925_ _18285_/Q _18284_/Q _12925_/C vssd1 vssd1 vccd1 vccd1 _12926_/C sky130_fd_sc_hd__and3_1
X_19481_ _19481_/CLK _19481_/D vssd1 vssd1 vccd1 vccd1 _19481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16097__S _16097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16693_ _16693_/A vssd1 vssd1 vccd1 vccd1 _16693_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18432_ _18818_/CLK _18432_/D vssd1 vssd1 vccd1 vccd1 _18432_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_61_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15644_ _15644_/A vssd1 vssd1 vccd1 vccd1 _18839_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _12897_/A _12863_/C vssd1 vssd1 vccd1 vccd1 _12856_/Y sky130_fd_sc_hd__nor2_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _19082_/CLK _18363_/D vssd1 vssd1 vccd1 vccd1 _18363_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _11733_/B _11740_/A _11806_/Y _11970_/A vssd1 vssd1 vccd1 vccd1 _11808_/B
+ sky130_fd_sc_hd__a31o_1
X_15575_ _18811_/Q _15574_/X _15584_/S vssd1 vssd1 vccd1 vccd1 _15576_/A sky130_fd_sc_hd__mux2_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _18534_/Q _18528_/Q _18527_/Q _18526_/Q vssd1 vssd1 vccd1 vccd1 _12789_/C
+ sky130_fd_sc_hd__or4b_1
XFILLER_15_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _17314_/A vssd1 vssd1 vccd1 vccd1 _19530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14526_ _16212_/B _14526_/B vssd1 vssd1 vccd1 vccd1 _14526_/Y sky130_fd_sc_hd__nand2_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18294_ _18298_/CLK _18294_/D vssd1 vssd1 vccd1 vccd1 _18294_/Q sky130_fd_sc_hd__dfxtp_2
X_11738_ _11738_/A vssd1 vssd1 vccd1 vccd1 _11738_/Y sky130_fd_sc_hd__inv_2
X_17245_ _19500_/Q _17244_/X _17245_/S vssd1 vssd1 vccd1 vccd1 _17246_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14457_ _18500_/Q _11984_/A _14465_/S vssd1 vssd1 vccd1 vccd1 _14458_/A sky130_fd_sc_hd__mux2_1
X_11669_ _12017_/B vssd1 vssd1 vccd1 vccd1 _12191_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13408_ _12850_/B _12582_/A _12584_/A _19853_/Q vssd1 vssd1 vccd1 vccd1 _13408_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_162_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17176_ _19479_/Q _17174_/X _17189_/S vssd1 vssd1 vccd1 vccd1 _17177_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14751__A2 _14703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14388_ _14388_/A vssd1 vssd1 vccd1 vccd1 _18474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16127_ _16127_/A vssd1 vssd1 vccd1 vccd1 _19042_/D sky130_fd_sc_hd__clkbuf_1
X_13339_ _19681_/Q _12737_/X _15242_/D _18405_/Q vssd1 vssd1 vccd1 vccd1 _13339_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16058_ _16768_/A vssd1 vssd1 vccd1 vccd1 _16058_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15009_ _16825_/A vssd1 vssd1 vccd1 vccd1 _15009_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15176__S _15185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09174__S _09190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19817_ _19818_/CLK _19817_/D vssd1 vssd1 vccd1 vccd1 _19817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19748_ _19759_/CLK _19748_/D vssd1 vssd1 vccd1 vccd1 _19748_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_110_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17205__A1 _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09501_ _09501_/A _09501_/B vssd1 vssd1 vccd1 vccd1 _09501_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19679_ _19682_/CLK _19679_/D vssd1 vssd1 vccd1 vccd1 _19679_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_38_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11733__A _11776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09432_ _18457_/Q _09309_/X _09396_/X _09431_/X vssd1 vssd1 vccd1 vccd1 _12505_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_53_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09363_ _09826_/A vssd1 vssd1 vccd1 vccd1 _09364_/A sky130_fd_sc_hd__buf_2
XANTENNA__10349__A _10349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16735__S _16735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11392__A_N _11722_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09294_ _18574_/Q _09255_/A _09291_/X _09293_/Y _18420_/Q vssd1 vssd1 vccd1 vccd1
+ _09303_/B sky130_fd_sc_hd__o221a_1
XFILLER_32_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16036__A _16135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_3_0_clock_A clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10439__S0 _11112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17566__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput150 _17884_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[15] sky130_fd_sc_hd__buf_2
XFILLER_82_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput161 _12322_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[25] sky130_fd_sc_hd__buf_2
XFILLER_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput172 _17866_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[6] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_30_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10611__S0 _10353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14258__A1 _12290_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12269__A0 _12265_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11167__S1 _10306_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10971_ _10873_/A _10966_/X _10970_/X _10827_/X vssd1 vssd1 vccd1 vccd1 _10971_/Y
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__09685__A1 _09402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12739__A _18290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12710_ _19803_/Q _12518_/X _12522_/X _18314_/Q _12709_/X vssd1 vssd1 vccd1 vccd1
+ _12711_/B sky130_fd_sc_hd__a221o_2
XFILLER_44_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13690_ _13688_/X _13689_/X _13758_/S vssd1 vssd1 vccd1 vccd1 _13690_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_3_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19610_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12458__B _12466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12641_ _12641_/A vssd1 vssd1 vccd1 vccd1 _13123_/A sky130_fd_sc_hd__buf_2
XFILLER_169_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13233__A2 _13230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15360_ _18729_/Q _15165_/X _15362_/S vssd1 vssd1 vccd1 vccd1 _15361_/A sky130_fd_sc_hd__mux2_1
X_12572_ _12572_/A vssd1 vssd1 vccd1 vccd1 _18340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17904__C1 _12802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14311_ _13979_/X _14312_/B _14309_/X _14310_/X vssd1 vssd1 vccd1 vccd1 _14311_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_168_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10452__C1 _10496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11523_ _12495_/A _13584_/A _13570_/D _11522_/X _11366_/A vssd1 vssd1 vccd1 vccd1
+ _11526_/B sky130_fd_sc_hd__a2111o_1
X_15291_ _15337_/S vssd1 vssd1 vccd1 vccd1 _15300_/S sky130_fd_sc_hd__buf_4
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17030_ _19419_/Q _16693_/X _17036_/S vssd1 vssd1 vccd1 vccd1 _17031_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14242_ _14312_/A _14237_/Y _14241_/Y _13864_/A vssd1 vssd1 vccd1 vccd1 _14242_/X
+ sky130_fd_sc_hd__o211a_1
X_11454_ _11458_/A vssd1 vssd1 vccd1 vccd1 _14426_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10405_ _10442_/A _10405_/B vssd1 vssd1 vccd1 vccd1 _10405_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14173_ _14173_/A vssd1 vssd1 vccd1 vccd1 _15123_/A sky130_fd_sc_hd__buf_4
X_11385_ _18424_/Q _11384_/Y _18425_/Q vssd1 vssd1 vccd1 vccd1 _11385_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_139_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13124_ _13428_/B vssd1 vssd1 vccd1 vccd1 _13205_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09783__A _09783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10336_ _19516_/Q _19130_/Q _19580_/Q _18736_/Q _10125_/A _09723_/A vssd1 vssd1 vccd1
+ vccd1 _10337_/B sky130_fd_sc_hd__mux4_1
XFILLER_140_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18981_ _18982_/CLK _18981_/D vssd1 vssd1 vccd1 vccd1 _18981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11818__A _19665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17932_ _17934_/B _17934_/C _17931_/Y vssd1 vssd1 vccd1 vccd1 _19762_/D sky130_fd_sc_hd__o21a_1
X_13055_ _13055_/A _18329_/Q _13055_/C vssd1 vssd1 vccd1 vccd1 _13056_/C sky130_fd_sc_hd__and3_1
XFILLER_140_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _19645_/Q _19062_/Q _19099_/Q _18705_/Q _11156_/S _09145_/A vssd1 vssd1 vccd1
+ vccd1 _10267_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12006_ _12481_/A _12004_/X _12126_/A vssd1 vssd1 vccd1 vccd1 _12008_/A sky130_fd_sc_hd__mux2_4
XFILLER_87_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17863_ _17863_/A vssd1 vssd1 vccd1 vccd1 _19732_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10602__S0 _10605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10198_ _19260_/Q _19031_/Q _18962_/Q _19356_/Q _10094_/A _09978_/A vssd1 vssd1 vccd1
+ vccd1 _10199_/B sky130_fd_sc_hd__mux4_1
XFILLER_121_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19602_ _19636_/CLK _19602_/D vssd1 vssd1 vccd1 vccd1 _19602_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15724__S _15730_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16814_ _16813_/X _19328_/Q _16823_/S vssd1 vssd1 vccd1 vccd1 _16815_/A sky130_fd_sc_hd__mux2_1
X_17794_ _15152_/X _19700_/Q _17794_/S vssd1 vssd1 vccd1 vccd1 _17795_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17199__A0 _19486_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16745_ _16826_/A vssd1 vssd1 vccd1 vccd1 _16845_/S sky130_fd_sc_hd__buf_8
X_19533_ _19534_/CLK _19533_/D vssd1 vssd1 vccd1 vccd1 _19533_/Q sky130_fd_sc_hd__dfxtp_1
X_13957_ _13969_/S _14103_/B vssd1 vssd1 vccd1 vccd1 _13957_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09220__S0 _09190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12908_ _12997_/A _12908_/B vssd1 vssd1 vccd1 vccd1 _12908_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19464_ _19592_/CLK _19464_/D vssd1 vssd1 vccd1 vccd1 _19464_/Q sky130_fd_sc_hd__dfxtp_1
X_16676_ _16676_/A vssd1 vssd1 vccd1 vccd1 _19285_/D sky130_fd_sc_hd__clkbuf_1
X_13888_ _13771_/X _13775_/X _13888_/S vssd1 vssd1 vccd1 vccd1 _13888_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18415_ _19481_/CLK _18415_/D vssd1 vssd1 vccd1 vccd1 _18415_/Q sky130_fd_sc_hd__dfxtp_2
X_15627_ _15649_/A vssd1 vssd1 vccd1 vccd1 _15636_/S sky130_fd_sc_hd__buf_4
XFILLER_62_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12839_ _12840_/B _12840_/C _18262_/Q vssd1 vssd1 vccd1 vccd1 _12841_/B sky130_fd_sc_hd__a21oi_1
X_19395_ _19395_/CLK _19395_/D vssd1 vssd1 vccd1 vccd1 _19395_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18981__D _18981_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14421__A1 _18518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18346_ _19759_/CLK _18346_/D vssd1 vssd1 vccd1 vccd1 _18346_/Q sky130_fd_sc_hd__dfxtp_1
X_15558_ _16813_/A vssd1 vssd1 vccd1 vccd1 _15558_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09523__S1 _09587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14509_ _17862_/A _14509_/B vssd1 vssd1 vccd1 vccd1 _14510_/A sky130_fd_sc_hd__or2_1
X_18277_ _18401_/CLK _18277_/D vssd1 vssd1 vccd1 vccd1 _18277_/Q sky130_fd_sc_hd__dfxtp_1
X_15489_ _16503_/A _15592_/B vssd1 vssd1 vccd1 vccd1 _15571_/A sky130_fd_sc_hd__nor2_2
XFILLER_163_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17228_ _17228_/A vssd1 vssd1 vccd1 vccd1 _19494_/D sky130_fd_sc_hd__clkbuf_1
Xinput30 io_dbus_rdata[7] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_4
Xinput41 io_ibus_inst[16] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__buf_2
Xinput52 io_ibus_inst[26] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__buf_2
XFILLER_156_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput63 io_ibus_inst[7] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17159_ _19474_/Q _17157_/X _17172_/S vssd1 vssd1 vccd1 vccd1 _17160_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16290__S _16296_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09981_ _09975_/Y _09977_/X _09980_/X _10022_/A vssd1 vssd1 vccd1 vccd1 _09981_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_170_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10632__A _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15634__S _15636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17415__A _17461_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12127__A1_N _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14660__A1 _14559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11463__A _11716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14660__B2 input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09415_ _09892_/A vssd1 vssd1 vccd1 vccd1 _09415_/X sky130_fd_sc_hd__buf_4
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12423__A0 _11202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ _10033_/S vssd1 vssd1 vccd1 vccd1 _09955_/A sky130_fd_sc_hd__buf_2
XANTENNA__09868__A _10029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ _09277_/A vssd1 vssd1 vccd1 vccd1 _09278_/A sky130_fd_sc_hd__buf_2
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10807__A _10807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17296__S _17302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11085__S0 _09447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11170_ _19625_/Q _19463_/Q _18909_/Q _18679_/Q _09692_/A _09704_/A vssd1 vssd1 vccd1
+ vccd1 _11171_/B sky130_fd_sc_hd__mux4_1
XFILLER_162_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14479__A1 _19748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_clock_A clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10121_ _19422_/Q _19198_/Q _19715_/Q _19166_/Q _10011_/S _09147_/A vssd1 vssd1 vccd1
+ vccd1 _10121_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13151__A1 _13139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ _19263_/Q _19034_/Q _18965_/Q _19359_/Q _09865_/A _10029_/A vssd1 vssd1 vccd1
+ vccd1 _10052_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14860_ _18439_/Q _14839_/S _14859_/X _14838_/A vssd1 vssd1 vccd1 vccd1 _14860_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13439__C1 _13401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13811_ _13811_/A vssd1 vssd1 vccd1 vccd1 _13811_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_35_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14791_ _16664_/A vssd1 vssd1 vccd1 vccd1 _16768_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input19_A io_dbus_rdata[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12469__A _12469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16530_ _19222_/Q _15526_/X _16536_/S vssd1 vssd1 vccd1 vccd1 _16531_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13742_ _13662_/X _13657_/X _13742_/S vssd1 vssd1 vccd1 vccd1 _13742_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_151_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19632_/CLK sky130_fd_sc_hd__clkbuf_16
X_10954_ _09926_/A _10944_/X _10953_/X _09305_/A _18429_/Q vssd1 vssd1 vccd1 vccd1
+ _12463_/A sky130_fd_sc_hd__a32o_4
XFILLER_44_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16461_ _16461_/A vssd1 vssd1 vccd1 vccd1 _19191_/D sky130_fd_sc_hd__clkbuf_1
X_13673_ _13670_/X _13672_/X _13747_/S vssd1 vssd1 vccd1 vccd1 _13673_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13206__A2 _12668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10885_ _10885_/A vssd1 vssd1 vccd1 vccd1 _10885_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18156__A _19839_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18200_ _19854_/Q _18200_/B vssd1 vssd1 vccd1 vccd1 _18201_/B sky130_fd_sc_hd__and2_1
XFILLER_25_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15412_ _16919_/A _15412_/B _15412_/C vssd1 vssd1 vccd1 vccd1 _16503_/B sky130_fd_sc_hd__or3_4
XFILLER_19_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12624_ _12624_/A vssd1 vssd1 vccd1 vccd1 _12703_/A sky130_fd_sc_hd__buf_2
XANTENNA__09778__A _09861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19180_ _19630_/CLK _19180_/D vssd1 vssd1 vccd1 vccd1 _19180_/Q sky130_fd_sc_hd__dfxtp_1
X_16392_ _16392_/A vssd1 vssd1 vccd1 vccd1 _19161_/D sky130_fd_sc_hd__clkbuf_1
X_18131_ _19830_/Q _18131_/B _18131_/C vssd1 vssd1 vccd1 vccd1 _18132_/C sky130_fd_sc_hd__and3_1
XANTENNA__10425__C1 _09459_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_166_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _18632_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11820__B _11820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15343_ _18721_/Q _15133_/X _15351_/S vssd1 vssd1 vccd1 vccd1 _15344_/A sky130_fd_sc_hd__mux2_1
X_12555_ _18419_/Q _12555_/B vssd1 vssd1 vccd1 vccd1 _12600_/A sky130_fd_sc_hd__and2b_2
XANTENNA__09830__A1 _09826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18062_ _18062_/A vssd1 vssd1 vccd1 vccd1 _18067_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11506_ _11506_/A _11506_/B vssd1 vssd1 vccd1 vccd1 _13529_/A sky130_fd_sc_hd__or2_2
XFILLER_7_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15274_ _18691_/Q _15146_/X _15278_/S vssd1 vssd1 vccd1 vccd1 _15275_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12486_ _12486_/A _12497_/B vssd1 vssd1 vccd1 vccd1 _12486_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12717__A1 _17774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17013_ _17013_/A vssd1 vssd1 vccd1 vccd1 _19411_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15719__S _15719_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14225_ _14059_/A _14227_/B _13975_/A _14224_/X vssd1 vssd1 vccd1 vccd1 _14225_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11437_ _18541_/Q _18540_/Q _12790_/A _18418_/Q vssd1 vssd1 vccd1 vccd1 _11438_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__12932__A _18288_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14156_ _13943_/A _14151_/Y _14155_/Y vssd1 vssd1 vccd1 vccd1 _14156_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_output87_A _12244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11368_ _11368_/A _11368_/B _11368_/C vssd1 vssd1 vccd1 vccd1 _11368_/X sky130_fd_sc_hd__and3_1
XFILLER_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13107_ _18347_/Q _12731_/A _13106_/X _13102_/X vssd1 vssd1 vccd1 vccd1 _18347_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _18768_/Q _18997_/Q _18928_/Q _19226_/Q _09692_/A _10306_/A vssd1 vssd1 vccd1
+ vccd1 _10320_/B sky130_fd_sc_hd__mux4_1
XFILLER_112_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18964_ _19584_/CLK _18964_/D vssd1 vssd1 vccd1 vccd1 _18964_/Q sky130_fd_sc_hd__dfxtp_1
X_14087_ _13918_/S _13890_/X _13899_/X vssd1 vssd1 vccd1 vccd1 _14087_/X sky130_fd_sc_hd__o21a_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15131__A2 _13873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _11299_/A _11664_/B vssd1 vssd1 vccd1 vccd1 _11575_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_104_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _18402_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13038_ _18324_/Q _13034_/C _13037_/Y vssd1 vssd1 vccd1 vccd1 _18324_/D sky130_fd_sc_hd__o21a_1
X_17915_ _19799_/Q _19801_/Q _19800_/Q _18036_/A vssd1 vssd1 vccd1 vccd1 _18046_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_112_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18895_ _19223_/CLK _18895_/D vssd1 vssd1 vccd1 vccd1 _18895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17846_ _17846_/A vssd1 vssd1 vccd1 vccd1 _19723_/D sky130_fd_sc_hd__clkbuf_1
X_17777_ _17779_/A _17777_/B vssd1 vssd1 vccd1 vccd1 _17778_/A sky130_fd_sc_hd__and2_2
X_14989_ input17/X _14960_/X _14925_/A vssd1 vssd1 vccd1 vccd1 _14994_/A sky130_fd_sc_hd__a21o_1
XFILLER_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_119_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _18578_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11456__A1 _14431_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19516_ _19612_/CLK _19516_/D vssd1 vssd1 vccd1 vccd1 _19516_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12653__B1 _12602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09744__S1 _09723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16728_ _16728_/A vssd1 vssd1 vccd1 vccd1 _16728_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11197__A2_N _09309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19447_ _19609_/CLK _19447_/D vssd1 vssd1 vccd1 vccd1 _19447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16659_ _19280_/Q _16657_/X _16671_/S vssd1 vssd1 vccd1 vccd1 _16660_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09200_ _11171_/A vssd1 vssd1 vccd1 vccd1 _10313_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09688__A _09688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19378_ _19540_/CLK _19378_/D vssd1 vssd1 vccd1 vccd1 _19378_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12956__A1 _18295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09131_ _10568_/A vssd1 vssd1 vccd1 vccd1 _10373_/A sky130_fd_sc_hd__clkbuf_4
X_18329_ _18329_/CLK _18329_/D vssd1 vssd1 vccd1 vccd1 _18329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10627__A _10875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13938__A _14274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13381__A1 _19686_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09680__S0 _09583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11458__A _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09964_ _19523_/Q _19137_/Q _19587_/Q _18743_/Q _09872_/S _09869_/A vssd1 vssd1 vccd1
+ vccd1 _09965_/B sky130_fd_sc_hd__mux4_1
XFILLER_104_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15122__A2 _15116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13133__A1 _19760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09895_ _09884_/X _09894_/X _09940_/A vssd1 vssd1 vccd1 vccd1 _09895_/X sky130_fd_sc_hd__mux2_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_14_0_clock_A clkbuf_3_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_83_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19687_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14708__S _14923_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09598__A _10389_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670_ _10813_/A vssd1 vssd1 vccd1 vccd1 _10670_/X sky130_fd_sc_hd__buf_2
XFILLER_139_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17335__A0 _16765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09329_ _09732_/A vssd1 vssd1 vccd1 vccd1 _11180_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__09812__A1 _09814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12340_ _18376_/Q _12341_/B vssd1 vssd1 vccd1 vccd1 _12340_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_98_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19791_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12271_ _11706_/X _12269_/X _12270_/X _12072_/X vssd1 vssd1 vccd1 vccd1 _12271_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12752__A _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14010_ _14003_/X _14006_/X _14007_/Y _14009_/X vssd1 vssd1 vccd1 vccd1 _14010_/Y
+ sky130_fd_sc_hd__o31ai_2
XFILLER_141_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11222_ _11222_/A _12500_/A vssd1 vssd1 vccd1 vccd1 _11222_/X sky130_fd_sc_hd__and2_1
XFILLER_107_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19452_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11153_ _11153_/A vssd1 vssd1 vccd1 vccd1 _11153_/X sky130_fd_sc_hd__buf_2
XFILLER_68_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10104_ _19520_/Q _19134_/Q _19584_/Q _18740_/Q _10094_/X _10103_/X vssd1 vssd1 vccd1
+ vccd1 _10105_/B sky130_fd_sc_hd__mux4_1
X_15961_ _16503_/B _17064_/B vssd1 vssd1 vccd1 vccd1 _16018_/A sky130_fd_sc_hd__or2_2
X_11084_ _11247_/A _11244_/A _11244_/B _11081_/Y _11083_/Y vssd1 vssd1 vccd1 vccd1
+ _11242_/C sky130_fd_sc_hd__o311ai_4
XFILLER_68_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15274__S _15278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10035_ _10042_/A _10030_/X _10032_/X _10034_/X vssd1 vssd1 vccd1 vccd1 _10035_/X
+ sky130_fd_sc_hd__o22a_1
X_17700_ _17700_/A vssd1 vssd1 vccd1 vccd1 _19676_/D sky130_fd_sc_hd__clkbuf_1
X_14912_ _18475_/Q _14912_/B vssd1 vssd1 vccd1 vccd1 _14932_/C sky130_fd_sc_hd__and2_1
X_15892_ _15892_/A vssd1 vssd1 vccd1 vccd1 _18949_/D sky130_fd_sc_hd__clkbuf_1
X_18680_ _19592_/CLK _18680_/D vssd1 vssd1 vccd1 vccd1 _18680_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_36_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19559_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17631_ _17631_/A vssd1 vssd1 vccd1 vccd1 _19664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14843_ _14861_/C _14841_/Y _14842_/X vssd1 vssd1 vccd1 vccd1 _14843_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_91_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17562_ _19640_/Q _16781_/A _17568_/S vssd1 vssd1 vccd1 vccd1 _17563_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14774_ _14772_/X _18591_/Q _14822_/S vssd1 vssd1 vccd1 vccd1 _14775_/A sky130_fd_sc_hd__mux2_1
X_11986_ _12408_/A vssd1 vssd1 vccd1 vccd1 _12294_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19301_ _19397_/CLK _19301_/D vssd1 vssd1 vccd1 vccd1 _19301_/Q sky130_fd_sc_hd__dfxtp_1
X_16513_ _16513_/A vssd1 vssd1 vccd1 vccd1 _19214_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13725_ _13893_/A vssd1 vssd1 vccd1 vccd1 _13950_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17493_ _17493_/A vssd1 vssd1 vccd1 vccd1 _19609_/D sky130_fd_sc_hd__clkbuf_1
X_10937_ _10933_/X _10935_/X _10936_/X _10701_/A _09407_/A vssd1 vssd1 vccd1 vccd1
+ _10944_/B sky130_fd_sc_hd__o221a_1
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_152_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19232_ _19620_/CLK _19232_/D vssd1 vssd1 vccd1 vccd1 _19232_/Q sky130_fd_sc_hd__dfxtp_1
X_16444_ _16501_/S vssd1 vssd1 vccd1 vccd1 _16453_/S sky130_fd_sc_hd__buf_2
X_13656_ _13629_/X _13652_/X _14103_/A vssd1 vssd1 vccd1 vccd1 _13656_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10868_ _10871_/A _10868_/B vssd1 vssd1 vccd1 vccd1 _10868_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12938__A1 _18289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12607_ _13222_/S vssd1 vssd1 vccd1 vccd1 _12669_/A sky130_fd_sc_hd__clkbuf_2
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19163_ _19712_/CLK _19163_/D vssd1 vssd1 vccd1 vccd1 _19163_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09301__A _18575_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16375_ _16375_/A vssd1 vssd1 vccd1 vccd1 _19153_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17326__A0 _16752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10447__A _10447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16833__S _16839_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13587_ _13587_/A _13587_/B _13587_/C vssd1 vssd1 vccd1 vccd1 _13720_/B sky130_fd_sc_hd__nand3_4
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10799_ _09409_/A _10787_/X _10792_/X _10798_/X vssd1 vssd1 vccd1 vccd1 _10799_/X
+ sky130_fd_sc_hd__a31o_2
X_18114_ _18114_/A _18119_/C vssd1 vssd1 vccd1 vccd1 _18114_/Y sky130_fd_sc_hd__nor2_1
X_15326_ _15326_/A vssd1 vssd1 vccd1 vccd1 _18714_/D sky130_fd_sc_hd__clkbuf_1
X_12538_ _12541_/B _12747_/C vssd1 vssd1 vccd1 vccd1 _12539_/A sky130_fd_sc_hd__nor2_1
X_19094_ _19640_/CLK _19094_/D vssd1 vssd1 vccd1 vccd1 _19094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18045_ _18077_/A _18045_/B _18045_/C vssd1 vssd1 vccd1 vccd1 _19800_/D sky130_fd_sc_hd__nor3_1
X_15257_ _15257_/A vssd1 vssd1 vccd1 vccd1 _18686_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12662__A _13130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12469_ _12469_/A _12469_/B vssd1 vssd1 vccd1 vccd1 _12469_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14208_ _12185_/X _14070_/A _14206_/X _14207_/Y vssd1 vssd1 vccd1 vccd1 _14208_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15188_ _15220_/A vssd1 vssd1 vccd1 vccd1 _15201_/S sky130_fd_sc_hd__buf_4
XFILLER_99_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14139_ _13937_/X _14138_/B _14040_/X vssd1 vssd1 vccd1 vccd1 _14139_/X sky130_fd_sc_hd__o21a_1
XFILLER_152_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18947_ _19633_/CLK _18947_/D vssd1 vssd1 vccd1 vccd1 _18947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14589__A _14589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09680_ _19430_/Q _19206_/Q _19723_/Q _19174_/Q _09583_/A _10451_/A vssd1 vssd1 vccd1
+ vccd1 _09680_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18878_ _19559_/CLK _18878_/D vssd1 vssd1 vccd1 vccd1 _18878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17829_ _17840_/A vssd1 vssd1 vccd1 vccd1 _17838_/S sky130_fd_sc_hd__buf_4
XFILLER_66_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12626__B1 _12742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16309__A _16355_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15213__A _16715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15040__A1 _13398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09114_ _11325_/C vssd1 vssd1 vccd1 vccd1 _11471_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11074__A2_N _12469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09653__S0 _09448_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09947_ _09947_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _09947_/X sky130_fd_sc_hd__or2_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11117__B1 _09393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14854__A1 _11542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10015__S1 _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ _09942_/A _09878_/B vssd1 vssd1 vccd1 vccd1 _09878_/Y sky130_fd_sc_hd__nor2_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10031__S _10033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11840_ _11840_/A vssd1 vssd1 vccd1 vccd1 _11948_/A sky130_fd_sc_hd__buf_2
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14946__B _14946_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _17762_/S _11770_/X _11997_/A vssd1 vssd1 vccd1 vccd1 _11771_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _18413_/Q _13423_/X _13512_/S vssd1 vssd1 vccd1 vccd1 _13511_/A sky130_fd_sc_hd__mux2_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15123__A _15123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10722_ _11065_/A vssd1 vssd1 vccd1 vccd1 _10797_/A sky130_fd_sc_hd__buf_2
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14490_ _18515_/Q _19753_/Q _14498_/S vssd1 vssd1 vccd1 vccd1 _14491_/A sky130_fd_sc_hd__mux2_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12466__B _12466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13441_ _13441_/A vssd1 vssd1 vccd1 vccd1 _18382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10653_ _18761_/Q _18990_/Q _18921_/Q _19219_/Q _10500_/A _09514_/A vssd1 vssd1 vccd1
+ vccd1 _10653_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11053__C1 _10797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16160_ _16160_/A vssd1 vssd1 vccd1 vccd1 _19054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13372_ _18329_/Q _13178_/X _12753_/A _19786_/Q vssd1 vssd1 vccd1 vccd1 _13372_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10584_ _10580_/X _10582_/X _10583_/X _10591_/A _10219_/A vssd1 vssd1 vccd1 vccd1
+ _10589_/B sky130_fd_sc_hd__o221a_1
XFILLER_155_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15111_ _15111_/A vssd1 vssd1 vccd1 vccd1 _15111_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12323_ _12323_/A vssd1 vssd1 vccd1 vccd1 _12419_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__13578__A _13578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16091_ _16090_/X _19031_/Q _16097_/S vssd1 vssd1 vccd1 vccd1 _16092_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12482__A _12482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15042_ _14999_/X _15036_/X _15039_/Y _15041_/X vssd1 vssd1 vccd1 vccd1 _16731_/A
+ sky130_fd_sc_hd__a22o_4
X_12254_ _13523_/B _12344_/A _12173_/Y vssd1 vssd1 vccd1 vccd1 _12254_/X sky130_fd_sc_hd__a21o_1
XFILLER_154_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12553__C1 _12552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11205_ _11205_/A _12505_/A vssd1 vssd1 vccd1 vccd1 _11205_/Y sky130_fd_sc_hd__nand2_1
X_19850_ _19851_/CLK _19850_/D vssd1 vssd1 vccd1 vccd1 _19850_/Q sky130_fd_sc_hd__dfxtp_2
X_12185_ _12185_/A _12185_/B vssd1 vssd1 vccd1 vccd1 _12185_/X sky130_fd_sc_hd__xor2_4
XANTENNA__10254__S1 _09697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15098__A1 _18624_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11529__C _13529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18801_ _19642_/CLK _18801_/D vssd1 vssd1 vccd1 vccd1 _18801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11136_ _11262_/A _11262_/B _11135_/X _10413_/A vssd1 vssd1 vccd1 vccd1 _11235_/C
+ sky130_fd_sc_hd__a211o_1
X_19781_ _19861_/CLK _19781_/D vssd1 vssd1 vccd1 vccd1 _19781_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10099__B_N _10098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16993_ _17049_/A vssd1 vssd1 vccd1 vccd1 _17062_/S sky130_fd_sc_hd__buf_6
X_18732_ _19640_/CLK _18732_/D vssd1 vssd1 vccd1 vccd1 _18732_/Q sky130_fd_sc_hd__dfxtp_1
X_15944_ _15044_/X _18973_/Q _15946_/S vssd1 vssd1 vccd1 vccd1 _15945_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11067_ _10774_/X _11060_/X _11062_/X _11066_/X _09390_/A vssd1 vssd1 vccd1 vccd1
+ _11067_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10018_ _10007_/X _10009_/X _10013_/X _10017_/X _09135_/A vssd1 vssd1 vccd1 vccd1
+ _10018_/X sky130_fd_sc_hd__a311o_1
XFILLER_92_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18663_ _19609_/CLK _18663_/D vssd1 vssd1 vccd1 vccd1 _18663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15875_ _15875_/A vssd1 vssd1 vccd1 vccd1 _18942_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15732__S _15734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17614_ _17707_/A vssd1 vssd1 vccd1 vccd1 _17625_/S sky130_fd_sc_hd__clkbuf_2
X_14826_ _18436_/Q _14839_/S _14824_/X _14838_/A vssd1 vssd1 vccd1 vccd1 _14826_/X
+ sky130_fd_sc_hd__o211a_1
X_18594_ _19704_/CLK _18594_/D vssd1 vssd1 vccd1 vccd1 _18594_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15270__A1 _15133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17545_ _17545_/A vssd1 vssd1 vccd1 vccd1 _19632_/D sky130_fd_sc_hd__clkbuf_1
X_14757_ _10810_/X _13181_/B _14922_/S vssd1 vssd1 vccd1 vccd1 _14757_/X sky130_fd_sc_hd__mux2_1
X_11969_ _11969_/A vssd1 vssd1 vccd1 vccd1 _14089_/B sky130_fd_sc_hd__buf_2
XFILLER_63_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11561__A _11561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13708_ _13922_/A _13922_/B vssd1 vssd1 vccd1 vccd1 _14276_/A sky130_fd_sc_hd__or2_1
X_17476_ _17533_/S vssd1 vssd1 vccd1 vccd1 _17485_/S sky130_fd_sc_hd__buf_2
X_14688_ _14694_/A _14688_/B vssd1 vssd1 vccd1 vccd1 _14689_/A sky130_fd_sc_hd__and2_1
X_19215_ _19698_/CLK _19215_/D vssd1 vssd1 vccd1 vccd1 _19215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13639_ _13769_/S vssd1 vssd1 vccd1 vccd1 _13776_/S sky130_fd_sc_hd__clkbuf_2
X_16427_ _16427_/A vssd1 vssd1 vccd1 vccd1 _19177_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16563__S _16569_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10177__A _10177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11044__C1 _19695_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16358_ _16503_/A _16992_/B vssd1 vssd1 vccd1 vccd1 _16415_/A sky130_fd_sc_hd__nor2_2
X_19146_ _19660_/CLK _19146_/D vssd1 vssd1 vccd1 vccd1 _19146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10398__A1 _09315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14591__B _14591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15179__S _15185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15309_ _18707_/Q _15197_/X _15311_/S vssd1 vssd1 vccd1 vccd1 _15310_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16289_ _16289_/A vssd1 vssd1 vccd1 vccd1 _19115_/D sky130_fd_sc_hd__clkbuf_1
X_19077_ _19647_/CLK _19077_/D vssd1 vssd1 vccd1 vccd1 _19077_/Q sky130_fd_sc_hd__dfxtp_1
X_18028_ _19795_/Q _18025_/B _18027_/Y vssd1 vssd1 vccd1 vccd1 _19795_/D sky130_fd_sc_hd__o21a_1
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17394__S _17402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15907__S _15913_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10116__S _10153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15089__A1 _11696_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09801_ _09278_/X _09786_/X _09800_/X _09285_/X _18450_/Q vssd1 vssd1 vccd1 vccd1
+ _11148_/A sky130_fd_sc_hd__a32o_4
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09732_ _09732_/A vssd1 vssd1 vccd1 vccd1 _11185_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09206__A _19694_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ _10245_/A vssd1 vssd1 vccd1 vccd1 _10390_/A sky130_fd_sc_hd__buf_4
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17786__A0 _15133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10322__A1 _09689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16738__S _16741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09594_ _18615_/Q _19304_/Q _10185_/S vssd1 vssd1 vccd1 vccd1 _09595_/B sky130_fd_sc_hd__mux2_1
XFILLER_27_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15013__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__S0 _10131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12378__A2 _14289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13327__B2 _18371_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_100_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15817__S _15819_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15118__A _15125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10550__A _10622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13990_ _18432_/Q _11460_/X _13989_/X vssd1 vssd1 vccd1 vccd1 _18432_/D sky130_fd_sc_hd__o21a_1
XANTENNA__11105__A3 _11104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12941_ _18291_/Q _12946_/C vssd1 vssd1 vccd1 vccd1 _12943_/B sky130_fd_sc_hd__nor2_1
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15552__S _15552_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15660_ _18847_/Q _15586_/X _15662_/S vssd1 vssd1 vccd1 vccd1 _15661_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12872_ _12873_/B _12873_/C _18271_/Q vssd1 vssd1 vccd1 vccd1 _12874_/B sky130_fd_sc_hd__a21oi_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _11468_/B _14597_/X _14593_/X _14610_/Y vssd1 vssd1 vccd1 vccd1 _14612_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11823_ _18355_/Q _11823_/B vssd1 vssd1 vccd1 vccd1 _11823_/Y sky130_fd_sc_hd__nor2_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _15591_/A vssd1 vssd1 vccd1 vccd1 _18816_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10077__B1 _09996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _16758_/X _19537_/Q _17330_/S vssd1 vssd1 vccd1 vccd1 _17331_/A sky130_fd_sc_hd__mux2_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _18565_/Q _14526_/B _14541_/Y _14535_/X vssd1 vssd1 vccd1 vccd1 _18533_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _11792_/B _11754_/B _12411_/B vssd1 vssd1 vccd1 vccd1 _11754_/X sky130_fd_sc_hd__or3b_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_25_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10172__S0 _09344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17479__S _17485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10705_ _10705_/A vssd1 vssd1 vccd1 vccd1 _10705_/Y sky130_fd_sc_hd__inv_2
X_17261_ _19506_/Q _16657_/X _17269_/S vssd1 vssd1 vccd1 vccd1 _17262_/A sky130_fd_sc_hd__mux2_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _14473_/A vssd1 vssd1 vccd1 vccd1 _18507_/D sky130_fd_sc_hd__clkbuf_1
X_11685_ _11685_/A vssd1 vssd1 vccd1 vccd1 _11685_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__16383__S _16391_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16212_ _16212_/A _16212_/B _16212_/C _16212_/D vssd1 vssd1 vccd1 vccd1 _17783_/A
+ sky130_fd_sc_hd__and4_4
X_19000_ _19165_/CLK _19000_/D vssd1 vssd1 vccd1 vccd1 _19000_/Q sky130_fd_sc_hd__dfxtp_1
X_13424_ _18380_/Q _13438_/B vssd1 vssd1 vccd1 vccd1 _13424_/X sky130_fd_sc_hd__or2_1
XFILLER_174_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17192_ _17226_/A vssd1 vssd1 vccd1 vccd1 _17206_/S sky130_fd_sc_hd__clkbuf_2
X_10636_ _10764_/A _10636_/B vssd1 vssd1 vccd1 vccd1 _10636_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16143_ _16143_/A vssd1 vssd1 vccd1 vccd1 _19046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13355_ _13390_/A _18644_/Q vssd1 vssd1 vccd1 vccd1 _13355_/Y sky130_fd_sc_hd__nand2_1
X_10567_ _09454_/A _10564_/X _10566_/X _09459_/A vssd1 vssd1 vccd1 vccd1 _10568_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13318__A1 _12617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13101__A input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12306_ _09898_/A _18515_/Q _12444_/S vssd1 vssd1 vccd1 vccd1 _12307_/A sky130_fd_sc_hd__mux2_4
X_16074_ _16784_/A vssd1 vssd1 vccd1 vccd1 _16074_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13286_ _19483_/Q _13235_/X _13236_/X _13295_/A _13285_/X vssd1 vssd1 vccd1 vccd1
+ _13288_/A sky130_fd_sc_hd__a221o_1
X_10498_ _10498_/A _10498_/B vssd1 vssd1 vccd1 vccd1 _10498_/X sky130_fd_sc_hd__or2_1
X_15025_ input20/X _14960_/X _15000_/X vssd1 vssd1 vccd1 vccd1 _15025_/X sky130_fd_sc_hd__a21o_1
X_12237_ _12237_/A _12237_/B vssd1 vssd1 vccd1 vccd1 _12237_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19833_ _19833_/CLK _19833_/D vssd1 vssd1 vccd1 vccd1 _19833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12168_ _13316_/A _12169_/C _18369_/Q vssd1 vssd1 vccd1 vccd1 _12168_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_151_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14818__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11119_ _11119_/A _11119_/B vssd1 vssd1 vccd1 vccd1 _11119_/Y sky130_fd_sc_hd__nor2_1
X_19764_ _19861_/CLK _19764_/D vssd1 vssd1 vccd1 vccd1 _19764_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10460__A _10461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12099_ _18366_/Q vssd1 vssd1 vccd1 vccd1 _13312_/A sky130_fd_sc_hd__clkbuf_2
X_16976_ _16976_/A vssd1 vssd1 vccd1 vccd1 _19395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18715_ _19722_/CLK _18715_/D vssd1 vssd1 vccd1 vccd1 _18715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15927_ _14951_/X _18965_/Q _15935_/S vssd1 vssd1 vccd1 vccd1 _15928_/A sky130_fd_sc_hd__mux2_1
Xinput6 io_dbus_rdata[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_2
XANTENNA__16558__S _16558_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19695_ _19695_/CLK _19695_/D vssd1 vssd1 vccd1 vccd1 _19695_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__10304__A1 _19061_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14867__A _16787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15462__S _15470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18646_ _19727_/CLK _18646_/D vssd1 vssd1 vccd1 vccd1 _18646_/Q sky130_fd_sc_hd__dfxtp_1
X_15858_ _15858_/A vssd1 vssd1 vccd1 vccd1 _18934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15243__A1 _16212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14809_ _14808_/X _18594_/Q _14822_/S vssd1 vssd1 vccd1 vccd1 _14810_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18577_ _18618_/CLK _18577_/D vssd1 vssd1 vccd1 vccd1 _18577_/Q sky130_fd_sc_hd__dfxtp_1
X_15789_ _14986_/X _18904_/Q _15791_/S vssd1 vssd1 vccd1 vccd1 _15790_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17528_ _17528_/A vssd1 vssd1 vccd1 vccd1 _19625_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11722__C _11722_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17389__S _17389_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17459_ _16841_/X _19595_/Q _17461_/S vssd1 vssd1 vccd1 vccd1 _17460_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17940__B1 _13063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14754__A0 _14753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09696__A _09704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19129_ _19579_/CLK _19129_/D vssd1 vssd1 vccd1 vccd1 _19129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12418__A1_N _14587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18248__A1 _18247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11466__A _15095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09715_ _18843_/Q _19397_/Q _19559_/Q _18811_/Q _09545_/S _10080_/A vssd1 vssd1 vccd1
+ vccd1 _09715_/X sky130_fd_sc_hd__mux4_1
XANTENNA__15880__B _17391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09646_ _09642_/X _09644_/X _09645_/X _09649_/A _09689_/A vssd1 vssd1 vccd1 vccd1
+ _09646_/X sky130_fd_sc_hd__o221a_1
XFILLER_83_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _18782_/Q _19011_/Q _18942_/Q _19240_/Q _09344_/A _10331_/A vssd1 vssd1 vccd1
+ vccd1 _09578_/B sky130_fd_sc_hd__mux4_2
XANTENNA__16992__A _16992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17931__B1 _13063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14745__B1 _14744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11470_ _11470_/A _12344_/A _14431_/C vssd1 vssd1 vccd1 vccd1 _13579_/B sky130_fd_sc_hd__or3_1
XANTENNA__09847__S0 _09914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10421_ _19415_/Q _19191_/Q _19708_/Q _19159_/Q _11087_/S _09142_/A vssd1 vssd1 vccd1
+ vccd1 _10421_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13140_ _13171_/A _18620_/Q vssd1 vssd1 vccd1 vccd1 _13140_/Y sky130_fd_sc_hd__nand2_1
X_10352_ _10733_/S vssd1 vssd1 vccd1 vccd1 _10353_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_151_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13071_ _17948_/A _18110_/C vssd1 vssd1 vccd1 vccd1 _13071_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10209__S1 _10080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10283_ _19419_/Q _19195_/Q _19712_/Q _19163_/Q _10224_/X _09486_/X vssd1 vssd1 vccd1
+ vccd1 _10283_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12760__A _14431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ _12043_/A _11928_/X _12018_/X _12021_/Y vssd1 vssd1 vccd1 vccd1 _17880_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09545__S _09545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09924__B1 _09425_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input49_A io_ibus_inst[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17762__S _17762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16830_ _16829_/X _19333_/Q _16839_/S vssd1 vssd1 vccd1 vccd1 _16831_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10280__A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13973_ _14122_/S _13972_/Y _13706_/A vssd1 vssd1 vccd1 vccd1 _13973_/Y sky130_fd_sc_hd__a21oi_1
X_16761_ _16761_/A vssd1 vssd1 vccd1 vccd1 _16761_/X sky130_fd_sc_hd__buf_2
XFILLER_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18500_ _18623_/CLK _18500_/D vssd1 vssd1 vccd1 vccd1 _18500_/Q sky130_fd_sc_hd__dfxtp_2
X_12924_ _12930_/C _12930_/D _12923_/Y vssd1 vssd1 vccd1 vccd1 _18285_/D sky130_fd_sc_hd__o21a_1
X_15712_ _15712_/A vssd1 vssd1 vccd1 vccd1 _18869_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19480_ _19488_/CLK _19480_/D vssd1 vssd1 vccd1 vccd1 _19480_/Q sky130_fd_sc_hd__dfxtp_1
X_16692_ _16692_/A vssd1 vssd1 vccd1 vccd1 _19290_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10393__S0 _10230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18431_ _19691_/CLK _18431_/D vssd1 vssd1 vccd1 vccd1 _18431_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_62_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12855_ _12865_/D vssd1 vssd1 vccd1 vccd1 _12863_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15643_ _18839_/Q _15561_/X _15647_/S vssd1 vssd1 vccd1 vccd1 _15644_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17998__A _18033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11806_ _13939_/B vssd1 vssd1 vccd1 vccd1 _11806_/Y sky130_fd_sc_hd__inv_2
X_18362_ _18381_/CLK _18362_/D vssd1 vssd1 vccd1 vccd1 _18362_/Q sky130_fd_sc_hd__dfxtp_1
X_15574_ _16829_/A vssd1 vssd1 vccd1 vccd1 _15574_/X sky130_fd_sc_hd__buf_2
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _18551_/Q _18550_/Q _18541_/Q _18540_/Q vssd1 vssd1 vccd1 vccd1 _12789_/B
+ sky130_fd_sc_hd__or4_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14525_ _18528_/Q _14522_/X _14524_/Y _14514_/X vssd1 vssd1 vccd1 vccd1 _18528_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _19530_/Q _16734_/X _17313_/S vssd1 vssd1 vccd1 vccd1 _17314_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _18565_/Q _11371_/Y _11535_/A _11736_/X vssd1 vssd1 vccd1 vccd1 _11738_/A
+ sky130_fd_sc_hd__o211a_1
X_18293_ _18298_/CLK _18293_/D vssd1 vssd1 vccd1 vccd1 _18293_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17244_ _18457_/Q _17628_/S _15263_/B vssd1 vssd1 vccd1 vccd1 _17244_/X sky130_fd_sc_hd__a21o_1
X_14456_ _14502_/S vssd1 vssd1 vccd1 vccd1 _14465_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_128_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11668_ _12219_/S _11663_/Y _11665_/X _11667_/X _11979_/A vssd1 vssd1 vccd1 vccd1
+ _11668_/X sky130_fd_sc_hd__a311o_1
XFILLER_30_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12654__B _14946_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13407_ _13407_/A _13407_/B vssd1 vssd1 vccd1 vccd1 _13407_/X sky130_fd_sc_hd__or2_1
XFILLER_174_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17175_ _17245_/S vssd1 vssd1 vccd1 vccd1 _17189_/S sky130_fd_sc_hd__clkbuf_2
X_10619_ _10750_/A _10611_/X _10618_/X _09225_/A vssd1 vssd1 vccd1 vccd1 _10619_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14387_ _18474_/Q _18506_/Q _14395_/S vssd1 vssd1 vccd1 vccd1 _14388_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11599_ _11599_/A _11599_/B _11599_/C vssd1 vssd1 vccd1 vccd1 _11686_/B sky130_fd_sc_hd__and3_1
XFILLER_128_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11050__S _11050_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16126_ _16125_/X _19042_/Q _16129_/S vssd1 vssd1 vccd1 vccd1 _16127_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13338_ _18289_/Q _12638_/X _13119_/C _18372_/Q vssd1 vssd1 vccd1 vccd1 _13338_/X
+ sky130_fd_sc_hd__a22o_2
XANTENNA__17150__A1 _18429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15457__S _15459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16057_ _16057_/A vssd1 vssd1 vccd1 vccd1 _19020_/D sky130_fd_sc_hd__clkbuf_1
X_13269_ _13403_/A _18632_/Q vssd1 vssd1 vccd1 vccd1 _13269_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15008_ _16721_/A vssd1 vssd1 vccd1 vccd1 _16825_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19816_ _19822_/CLK _19816_/D vssd1 vssd1 vccd1 vccd1 _19816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19747_ _19755_/CLK _19747_/D vssd1 vssd1 vccd1 vccd1 _19747_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16288__S _16296_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12278__B2 _12497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16959_ _16959_/A vssd1 vssd1 vccd1 vccd1 _19387_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18069__A _18077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14597__A _18205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09500_ _18616_/Q _19305_/Q _10401_/A vssd1 vssd1 vccd1 vccd1 _09501_/B sky130_fd_sc_hd__mux2_1
XANTENNA__15192__S _15201_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19678_ _19680_/CLK _19678_/D vssd1 vssd1 vccd1 vccd1 _19678_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_64_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09431_ _09940_/A _09424_/X _09430_/X vssd1 vssd1 vccd1 vccd1 _09431_/X sky130_fd_sc_hd__a21o_1
XFILLER_53_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18629_ _18632_/CLK _18629_/D vssd1 vssd1 vccd1 vccd1 _18629_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11537__A_N _13570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15920__S _15924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09362_ _09810_/A vssd1 vssd1 vccd1 vccd1 _09826_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_162_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16716__A1 _16715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11253__A2 _12458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ _18576_/Q _15134_/A vssd1 vssd1 vccd1 vccd1 _09293_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14727__B1 _14726_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17847__S _17849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12202__A1 _18575_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10439__S1 _09602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10365__A _10365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13676__A _13845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15367__S _15373_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput140 _12469_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[7] sky130_fd_sc_hd__buf_2
XANTENNA__16052__A _16135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput151 _12103_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[16] sky130_fd_sc_hd__buf_2
XFILLER_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput162 _12343_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[26] sky130_fd_sc_hd__buf_2
Xoutput173 _17868_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[7] sky130_fd_sc_hd__buf_2
XFILLER_43_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17582__S _17590_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10611__S1 _10548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15455__A1 _15194_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10970_ _09169_/A _10967_/X _10969_/X _10973_/A vssd1 vssd1 vccd1 vccd1 _10970_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_56_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09629_ _09629_/A vssd1 vssd1 vccd1 vccd1 _10560_/S sky130_fd_sc_hd__buf_2
XFILLER_15_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12640_ _12640_/A vssd1 vssd1 vccd1 vccd1 _12641_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12571_ _12559_/X _12562_/X _13092_/S vssd1 vssd1 vccd1 vccd1 _12572_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12441__A1 _19758_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16707__A1 _16705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14310_ _14332_/A _14310_/B vssd1 vssd1 vccd1 vccd1 _14310_/X sky130_fd_sc_hd__or2_1
XFILLER_157_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11522_ _11522_/A _11522_/B _11549_/A vssd1 vssd1 vccd1 vccd1 _11522_/X sky130_fd_sc_hd__and3_1
XFILLER_11_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15290_ _15290_/A vssd1 vssd1 vccd1 vccd1 _18698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12474__B _12474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14241_ _14241_/A _14241_/B vssd1 vssd1 vccd1 vccd1 _14241_/Y sky130_fd_sc_hd__nand2_1
X_11453_ input72/X _14431_/A vssd1 vssd1 vccd1 vccd1 _11458_/A sky130_fd_sc_hd__nor2_2
X_10404_ _19515_/Q _19129_/Q _19579_/Q _18735_/Q _10224_/X _11111_/A vssd1 vssd1 vccd1
+ vccd1 _10405_/B sky130_fd_sc_hd__mux4_1
XFILLER_171_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14172_ _14328_/A _14172_/B vssd1 vssd1 vccd1 vccd1 _14172_/Y sky130_fd_sc_hd__nand2_1
X_11384_ _18426_/Q vssd1 vssd1 vccd1 vccd1 _11384_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13123_ _13123_/A vssd1 vssd1 vccd1 vccd1 _13123_/X sky130_fd_sc_hd__clkbuf_2
X_10335_ _09616_/X _10325_/Y _10327_/Y _09394_/A _10334_/X vssd1 vssd1 vccd1 vccd1
+ _10335_/X sky130_fd_sc_hd__o311a_2
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18980_ _18982_/CLK _18980_/D vssd1 vssd1 vccd1 vccd1 _18980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17931_ _17934_/B _17934_/C _13063_/X vssd1 vssd1 vccd1 vccd1 _17931_/Y sky130_fd_sc_hd__a21oi_1
X_13054_ _13055_/A _13055_/C _18329_/Q vssd1 vssd1 vccd1 vccd1 _13056_/B sky130_fd_sc_hd__a21oi_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10266_ _10270_/A _10266_/B vssd1 vssd1 vccd1 vccd1 _10266_/X sky130_fd_sc_hd__or2_1
XFILLER_30_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17492__S _17496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12005_ _12005_/A vssd1 vssd1 vccd1 vccd1 _12126_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17862_ _17862_/A _17862_/B vssd1 vssd1 vccd1 vccd1 _17863_/A sky130_fd_sc_hd__or2_1
XFILLER_121_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10602__S1 _10366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10197_ _10197_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _11230_/A sky130_fd_sc_hd__nor2_1
XANTENNA__15446__A1 _15181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19601_ _19601_/CLK _19601_/D vssd1 vssd1 vccd1 vccd1 _19601_/Q sky130_fd_sc_hd__dfxtp_1
X_16813_ _16813_/A vssd1 vssd1 vccd1 vccd1 _16813_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17793_ _17793_/A vssd1 vssd1 vccd1 vccd1 _19699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19532_ _19727_/CLK _19532_/D vssd1 vssd1 vccd1 vccd1 _19532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16744_ _16744_/A _17064_/B vssd1 vssd1 vccd1 vccd1 _16826_/A sky130_fd_sc_hd__or2_2
X_13956_ _13997_/S _13766_/X _13955_/X vssd1 vssd1 vccd1 vccd1 _14103_/B sky130_fd_sc_hd__o21ai_1
XFILLER_81_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09220__S1 _09149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12907_ _18281_/Q _12907_/B vssd1 vssd1 vccd1 vccd1 _12908_/B sky130_fd_sc_hd__and2_1
X_19463_ _19590_/CLK _19463_/D vssd1 vssd1 vccd1 vccd1 _19463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13887_ _13839_/S _13818_/B _13965_/S vssd1 vssd1 vccd1 vccd1 _13887_/Y sky130_fd_sc_hd__a21oi_1
X_16675_ _19285_/Q _16673_/X _16687_/S vssd1 vssd1 vccd1 vccd1 _16676_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16836__S _16839_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18414_ _19780_/CLK _18414_/D vssd1 vssd1 vccd1 vccd1 _18414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12838_ _12840_/B _12840_/C _12837_/Y vssd1 vssd1 vccd1 vccd1 _18261_/D sky130_fd_sc_hd__o21a_1
X_15626_ _15626_/A vssd1 vssd1 vccd1 vccd1 _18831_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19394_ _19556_/CLK _19394_/D vssd1 vssd1 vccd1 vccd1 _19394_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18345_ _18402_/CLK _18345_/D vssd1 vssd1 vccd1 vccd1 _18345_/Q sky130_fd_sc_hd__dfxtp_1
X_12769_ _18291_/Q _13404_/B vssd1 vssd1 vccd1 vccd1 _12769_/X sky130_fd_sc_hd__and2_1
X_15557_ _15557_/A vssd1 vssd1 vccd1 vccd1 _18805_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10884__S _10932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14508_ _11297_/B _18523_/Q _14516_/S vssd1 vssd1 vccd1 vccd1 _14509_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18276_ _18401_/CLK _18276_/D vssd1 vssd1 vccd1 vccd1 _18276_/Q sky130_fd_sc_hd__dfxtp_1
X_15488_ _16430_/A _16357_/B _16919_/C vssd1 vssd1 vccd1 vccd1 _15592_/B sky130_fd_sc_hd__or3b_4
XFILLER_30_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10994__A1 _10956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14185__A1 _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17227_ _19494_/Q _17225_/X _17239_/S vssd1 vssd1 vccd1 vccd1 _17228_/A sky130_fd_sc_hd__mux2_1
Xinput20 io_dbus_rdata[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_2
Xinput31 io_dbus_rdata[8] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_2
XANTENNA__16571__S _16573_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14439_ _18492_/Q _19730_/Q _14443_/S vssd1 vssd1 vccd1 vccd1 _14440_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput42 io_ibus_inst[17] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__buf_2
Xinput53 io_ibus_inst[27] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__buf_2
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput64 io_ibus_inst[8] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_1
X_17158_ _17245_/S vssd1 vssd1 vccd1 vccd1 _17172_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_171_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16109_ _16819_/A vssd1 vssd1 vccd1 vccd1 _16109_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09980_ _19265_/Q _19036_/Q _18967_/Q _19361_/Q _09782_/A _09979_/X vssd1 vssd1 vccd1
+ vccd1 _09980_/X sky130_fd_sc_hd__mux4_1
X_17089_ _16777_/X _19445_/Q _17097_/S vssd1 vssd1 vccd1 vccd1 _17090_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_147_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15437__A1 _15168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15216__A _16718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14120__A _14120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09214__A _09214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14660__A2 _12660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15650__S _15658_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09414_ _09414_/A vssd1 vssd1 vccd1 vccd1 _09892_/A sky130_fd_sc_hd__buf_2
XFILLER_41_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09345_ _10055_/S vssd1 vssd1 vccd1 vccd1 _10033_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_80_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10434__B1 _09459_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09276_ _09276_/A vssd1 vssd1 vccd1 vccd1 _09277_/A sky130_fd_sc_hd__buf_2
XFILLER_32_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10985__A1 _10548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17577__S _17579_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11085__S1 _09635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10823__A _10823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10120_ _10120_/A _10120_/B vssd1 vssd1 vccd1 vccd1 _10120_/X sky130_fd_sc_hd__or2_1
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13151__A2 _13149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ _10051_/A _12491_/C vssd1 vssd1 vccd1 vccd1 _11269_/B sky130_fd_sc_hd__or2b_1
XFILLER_88_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14100__A1 _11978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ _13810_/A vssd1 vssd1 vccd1 vccd1 _13810_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14790_ input30/X _14703_/A _14789_/X _14732_/X vssd1 vssd1 vccd1 vccd1 _16664_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_63_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13741_ _13659_/X _13681_/X _13741_/S vssd1 vssd1 vccd1 vccd1 _13741_/X sky130_fd_sc_hd__mux2_1
X_10953_ _10946_/X _10948_/X _10950_/X _10952_/X _09391_/A vssd1 vssd1 vccd1 vccd1
+ _10953_/X sky130_fd_sc_hd__a221o_1
XFILLER_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13672_ _12424_/A _13800_/B _13724_/B vssd1 vssd1 vccd1 vccd1 _13672_/X sky130_fd_sc_hd__mux2_1
X_16460_ _16074_/X _19191_/Q _16464_/S vssd1 vssd1 vccd1 vccd1 _16461_/A sky130_fd_sc_hd__mux2_1
X_10884_ _18851_/Q _19309_/Q _10932_/S vssd1 vssd1 vccd1 vccd1 _10885_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15061__C1 _14893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18156__B _19838_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12623_ _18286_/Q _13156_/A _12531_/Y _18337_/Q vssd1 vssd1 vccd1 vccd1 _12623_/X
+ sky130_fd_sc_hd__a22o_1
X_15411_ _15411_/A vssd1 vssd1 vccd1 vccd1 _18752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16391_ _19161_/Q _15535_/X _16391_/S vssd1 vssd1 vccd1 vccd1 _16392_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12485__A _12485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18130_ _18131_/B _18131_/C _19830_/Q vssd1 vssd1 vccd1 vccd1 _18132_/B sky130_fd_sc_hd__a21oi_1
XFILLER_129_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15342_ _15410_/S vssd1 vssd1 vccd1 vccd1 _15351_/S sky130_fd_sc_hd__clkbuf_4
X_12554_ _18635_/Q _12554_/B vssd1 vssd1 vccd1 vccd1 _12554_/X sky130_fd_sc_hd__or2_1
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11505_ _11665_/B _11664_/A _11664_/D _11512_/A vssd1 vssd1 vccd1 vccd1 _11506_/B
+ sky130_fd_sc_hd__or4_1
X_18061_ _18077_/A _18061_/B _18061_/C vssd1 vssd1 vccd1 vccd1 _19806_/D sky130_fd_sc_hd__nor3_1
X_15273_ _15273_/A vssd1 vssd1 vccd1 vccd1 _18690_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16391__S _16391_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12485_ _12485_/A _12497_/B vssd1 vssd1 vccd1 vccd1 _12485_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12178__A0 _10098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17012_ _19411_/Q _16667_/X _17014_/S vssd1 vssd1 vccd1 vccd1 _17013_/A sky130_fd_sc_hd__mux2_1
X_14224_ _14262_/A _14227_/A vssd1 vssd1 vccd1 vccd1 _14224_/X sky130_fd_sc_hd__and2_1
X_11436_ _18539_/Q _18538_/Q _18537_/Q vssd1 vssd1 vccd1 vccd1 _12790_/A sky130_fd_sc_hd__or3_1
XFILLER_137_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14155_ _14155_/A _14155_/B vssd1 vssd1 vccd1 vccd1 _14155_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11367_ _11580_/C _13579_/A _11367_/C _11367_/D vssd1 vssd1 vccd1 vccd1 _11593_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_99_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15667__A1 _15487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13106_ input71/X _13106_/B vssd1 vssd1 vccd1 vccd1 _13106_/X sky130_fd_sc_hd__or2_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _19418_/Q _19194_/Q _19711_/Q _19162_/Q _09701_/S _10306_/X vssd1 vssd1 vccd1
+ vccd1 _10318_/X sky130_fd_sc_hd__mux4_1
X_14086_ _13898_/X _14085_/X _14086_/S vssd1 vssd1 vccd1 vccd1 _14086_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13678__A0 _13623_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18963_ _19165_/CLK _18963_/D vssd1 vssd1 vccd1 vccd1 _18963_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _14513_/A _11298_/B vssd1 vssd1 vccd1 vccd1 _11664_/B sky130_fd_sc_hd__nand2_1
XFILLER_140_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _13049_/A _13045_/C vssd1 vssd1 vccd1 vccd1 _13037_/Y sky130_fd_sc_hd__nor2_1
X_17914_ _19797_/Q _19796_/Q _19798_/Q _18026_/A vssd1 vssd1 vccd1 vccd1 _18036_/A
+ sky130_fd_sc_hd__and4_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10249_ _11119_/A _10246_/X _10248_/X vssd1 vssd1 vccd1 vccd1 _10249_/Y sky130_fd_sc_hd__o21ai_1
X_18894_ _19513_/CLK _18894_/D vssd1 vssd1 vccd1 vccd1 _18894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17845_ _15226_/X _19723_/Q _17849_/S vssd1 vssd1 vccd1 vccd1 _17846_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17776_ _17776_/A vssd1 vssd1 vccd1 vccd1 _19692_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14988_ _14988_/A vssd1 vssd1 vccd1 vccd1 _18609_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19515_ _19643_/CLK _19515_/D vssd1 vssd1 vccd1 vccd1 _19515_/Q sky130_fd_sc_hd__dfxtp_1
X_16727_ _16727_/A vssd1 vssd1 vccd1 vccd1 _19301_/D sky130_fd_sc_hd__clkbuf_1
X_13939_ _14178_/A _13939_/B vssd1 vssd1 vccd1 vccd1 _13939_/X sky130_fd_sc_hd__or2_1
XFILLER_34_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15470__S _15470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09969__A _09969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19446_ _19608_/CLK _19446_/D vssd1 vssd1 vccd1 vccd1 _19446_/Q sky130_fd_sc_hd__dfxtp_1
X_16658_ _16741_/S vssd1 vssd1 vccd1 vccd1 _16671_/S sky130_fd_sc_hd__buf_2
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15609_ _15609_/A vssd1 vssd1 vccd1 vccd1 _18823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19377_ _19539_/CLK _19377_/D vssd1 vssd1 vccd1 vccd1 _19377_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09688__B _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16589_ _19250_/Q vssd1 vssd1 vccd1 vccd1 _16590_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_73_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09130_ _10823_/A vssd1 vssd1 vccd1 vccd1 _10568_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18328_ _18330_/CLK _18328_/D vssd1 vssd1 vccd1 vccd1 _18328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18259_ _19855_/CLK _18259_/D vssd1 vssd1 vccd1 vccd1 _18259_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18082__A _18170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11916__A0 _10554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_2_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19513_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09680__S1 _10451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09963_ _09892_/X _09958_/X _09960_/X _09962_/X _09940_/A vssd1 vssd1 vccd1 vccd1
+ _09963_/X sky130_fd_sc_hd__a221o_2
XANTENNA__15645__S _15647_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14330__A1 _18456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09894_ _09415_/X _09886_/Y _09888_/Y _09890_/Y _09893_/Y vssd1 vssd1 vccd1 vccd1
+ _09894_/X sky130_fd_sc_hd__o32a_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10789__S _10886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15380__S _15384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11921__B _13614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09328_ _10288_/A vssd1 vssd1 vccd1 vccd1 _09732_/A sky130_fd_sc_hd__buf_2
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14149__A1 _18441_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09259_ _18572_/Q _14716_/A vssd1 vssd1 vccd1 vccd1 _09259_/X sky130_fd_sc_hd__and2_1
XFILLER_167_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16505__A _16573_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17100__S _17108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _19682_/Q _12390_/B vssd1 vssd1 vccd1 vccd1 _12270_/X sky130_fd_sc_hd__or2_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11221_ _11225_/B _11225_/C _11152_/D _09899_/Y vssd1 vssd1 vccd1 vccd1 _11221_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12175__A3 _14192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11152_ _11225_/B _11225_/C _11152_/C _11152_/D vssd1 vssd1 vccd1 vccd1 _11152_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_161_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10103_ _10103_/A vssd1 vssd1 vccd1 vccd1 _10103_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__14321__A1 _11602_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15960_ _16212_/A _16212_/B _15960_/C vssd1 vssd1 vccd1 vccd1 _17064_/B sky130_fd_sc_hd__or3_4
X_11083_ _11083_/A vssd1 vssd1 vccd1 vccd1 _11083_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10569__S0 _10466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input31_A io_dbus_rdata[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _09881_/A _10033_/X _10068_/A vssd1 vssd1 vccd1 vccd1 _10034_/X sky130_fd_sc_hd__a21o_1
X_14911_ _18443_/Q _12594_/B _15071_/S vssd1 vssd1 vccd1 vccd1 _14911_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15891_ _14761_/X _18949_/Q _15891_/S vssd1 vssd1 vccd1 vccd1 _15892_/A sky130_fd_sc_hd__mux2_1
X_17630_ _19664_/Q _17628_/X _17653_/S vssd1 vssd1 vccd1 vccd1 _17631_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14842_ _14842_/A vssd1 vssd1 vccd1 vccd1 _14842_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17561_ _17561_/A vssd1 vssd1 vccd1 vccd1 _19639_/D sky130_fd_sc_hd__clkbuf_1
X_11985_ _11985_/A _12067_/D vssd1 vssd1 vccd1 vccd1 _11985_/Y sky130_fd_sc_hd__nor2_1
X_14773_ _15077_/S vssd1 vssd1 vccd1 vccd1 _14822_/S sky130_fd_sc_hd__clkbuf_4
X_19300_ _19622_/CLK _19300_/D vssd1 vssd1 vccd1 vccd1 _19300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16512_ _19214_/Q _15500_/X _16514_/S vssd1 vssd1 vccd1 vccd1 _16513_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10936_ _19246_/Q _19017_/Q _18948_/Q _19342_/Q _10886_/S _09352_/A vssd1 vssd1 vccd1
+ vccd1 _10936_/X sky130_fd_sc_hd__mux4_2
X_13724_ _13729_/B _13724_/B vssd1 vssd1 vccd1 vccd1 _13893_/A sky130_fd_sc_hd__and2_1
XFILLER_56_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17492_ _19609_/Q _16680_/X _17496_/S vssd1 vssd1 vccd1 vccd1 _17493_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19231_ _19553_/CLK _19231_/D vssd1 vssd1 vccd1 vccd1 _19231_/Q sky130_fd_sc_hd__dfxtp_1
X_16443_ _16443_/A vssd1 vssd1 vccd1 vccd1 _19183_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13655_ _13995_/S vssd1 vssd1 vccd1 vccd1 _14103_/A sky130_fd_sc_hd__clkbuf_2
X_10867_ _19408_/Q _19184_/Q _19701_/Q _19152_/Q _10664_/S _10365_/A vssd1 vssd1 vccd1
+ vccd1 _10868_/B sky130_fd_sc_hd__mux4_1
XFILLER_158_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12606_ _12606_/A vssd1 vssd1 vccd1 vccd1 _13404_/B sky130_fd_sc_hd__clkbuf_2
X_19162_ _19551_/CLK _19162_/D vssd1 vssd1 vccd1 vccd1 _19162_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16374_ _19153_/Q _15510_/X _16380_/S vssd1 vssd1 vccd1 vccd1 _16375_/A sky130_fd_sc_hd__mux2_1
X_13586_ _11355_/Y _11343_/X _11356_/Y _13585_/X _11366_/B vssd1 vssd1 vccd1 vccd1
+ _13587_/C sky130_fd_sc_hd__a311oi_4
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10798_ _10793_/X _10795_/X _10797_/X _10944_/A vssd1 vssd1 vccd1 vccd1 _10798_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_169_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18113_ _18122_/D vssd1 vssd1 vccd1 vccd1 _18119_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_12537_ _12686_/A _12537_/B vssd1 vssd1 vccd1 vccd1 _12541_/B sky130_fd_sc_hd__or2_2
X_15325_ _18714_/Q _15219_/X _15333_/S vssd1 vssd1 vccd1 vccd1 _15326_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19093_ _19706_/CLK _19093_/D vssd1 vssd1 vccd1 vccd1 _19093_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13348__C1 _13317_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17010__S _17014_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18044_ _18043_/A _18043_/C _19800_/Q vssd1 vssd1 vccd1 vccd1 _18045_/C sky130_fd_sc_hd__a21oi_1
X_15256_ _18686_/Q _15255_/X _15260_/S vssd1 vssd1 vccd1 vccd1 _15257_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12468_ _12468_/A _12469_/B vssd1 vssd1 vccd1 vccd1 _12468_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11419_ _12519_/A _12520_/A _11419_/C vssd1 vssd1 vccd1 vccd1 _12603_/A sky130_fd_sc_hd__nor3_4
XANTENNA__11559__A _16212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14207_ _13832_/A _14073_/Y _14012_/X vssd1 vssd1 vccd1 vccd1 _14207_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_160_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15187_ _16689_/A vssd1 vssd1 vccd1 vccd1 _15187_/X sky130_fd_sc_hd__buf_2
XFILLER_153_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12399_ _14310_/B _12399_/B vssd1 vssd1 vccd1 vccd1 _12403_/A sky130_fd_sc_hd__xor2_1
XANTENNA__12571__A0 _12559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14138_ _14140_/B _14138_/B vssd1 vssd1 vccd1 vccd1 _14142_/B sky130_fd_sc_hd__and2_1
XFILLER_153_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18946_ _19699_/CLK _18946_/D vssd1 vssd1 vccd1 vccd1 _18946_/Q sky130_fd_sc_hd__dfxtp_1
X_14069_ _18436_/Q _11460_/X _14068_/X vssd1 vssd1 vccd1 vccd1 _18436_/D sky130_fd_sc_hd__o21a_1
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18877_ _19559_/CLK _18877_/D vssd1 vssd1 vccd1 vccd1 _18877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17828_ _17828_/A vssd1 vssd1 vccd1 vccd1 _19715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12626__A1 _19678_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17759_ _17730_/X _13399_/X _17625_/S vssd1 vssd1 vccd1 vccd1 _17759_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__16296__S _16296_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14809__S _14822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18077__A _18077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19429_ _19591_/CLK _19429_/D vssd1 vssd1 vccd1 vccd1 _19429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09113_ _09113_/A _09113_/B vssd1 vssd1 vccd1 vccd1 _13570_/B sky130_fd_sc_hd__nor2_8
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12853__A _18170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10373__A _10373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_150_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19598_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09653__S1 _10349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09946_ _19620_/Q _19458_/Q _18904_/Q _18674_/Q _09955_/A _09881_/A vssd1 vssd1 vccd1
+ vccd1 _09947_/B sky130_fd_sc_hd__mux4_1
XANTENNA__11117__A1 _10219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_165_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19634_/CLK sky130_fd_sc_hd__clkbuf_16
X_09877_ _18778_/Q _19007_/Q _18938_/Q _19236_/Q _09803_/X _09810_/X vssd1 vssd1 vccd1
+ vccd1 _09878_/B sky130_fd_sc_hd__mux4_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17590__S _17590_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11932__A _11984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14946__C _14946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _18354_/Q _11758_/X _11768_/Y _11769_/X vssd1 vssd1 vccd1 vccd1 _11770_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13290__B2 _18247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11651__B _13665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10721_ _10946_/A _10721_/B vssd1 vssd1 vccd1 vccd1 _10721_/X sky130_fd_sc_hd__or2_1
XANTENNA__09402__A _09402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10548__A _10548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _13112_/A _18382_/Q _13440_/S vssd1 vssd1 vccd1 vccd1 _13441_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10652_ _09662_/A _10649_/Y _10651_/Y _10764_/A vssd1 vssd1 vccd1 vccd1 _10652_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_103_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _18401_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_142_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13371_ _12840_/B _12604_/X _12749_/X _19818_/Q vssd1 vssd1 vccd1 vccd1 _13371_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10982__S _10982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14790__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10583_ _19252_/Q _19023_/Q _18954_/Q _19348_/Q _10581_/S _09662_/A vssd1 vssd1 vccd1
+ vccd1 _10583_/X sky130_fd_sc_hd__mux4_1
XANTENNA__14790__B2 _14732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12763__A _14519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12322_ _12318_/Y _12321_/X _19753_/Q _12002_/X vssd1 vssd1 vccd1 vccd1 _12322_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_15110_ _18633_/Q _15109_/X _15104_/X _10412_/A vssd1 vssd1 vccd1 vccd1 _18633_/D
+ sky130_fd_sc_hd__a22o_1
X_16090_ _16800_/A vssd1 vssd1 vccd1 vccd1 _16090_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15041_ _14744_/X _15040_/X _14842_/X vssd1 vssd1 vccd1 vccd1 _15041_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12253_ _12246_/A _12116_/X _12249_/X _12252_/Y vssd1 vssd1 vccd1 vccd1 _17898_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__14542__A1 _18565_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_118_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _18618_/CLK sky130_fd_sc_hd__clkbuf_16
X_11204_ _11220_/A _11220_/B _11249_/A vssd1 vssd1 vccd1 vccd1 _11204_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_134_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12184_ _12141_/A _12141_/B _12163_/A _12183_/X vssd1 vssd1 vccd1 vccd1 _12185_/B
+ sky130_fd_sc_hd__a31o_2
XANTENNA__15098__A2 _13566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18800_ _19549_/CLK _18800_/D vssd1 vssd1 vccd1 vccd1 _18800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17066__A _17134_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11135_ _11135_/A _12483_/A vssd1 vssd1 vccd1 vccd1 _11135_/X sky130_fd_sc_hd__and2_1
X_19780_ _19780_/CLK _19780_/D vssd1 vssd1 vccd1 vccd1 _19780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16992_ _16992_/A _16992_/B vssd1 vssd1 vccd1 vccd1 _17049_/A sky130_fd_sc_hd__nor2_4
XFILLER_62_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18731_ _19639_/CLK _18731_/D vssd1 vssd1 vccd1 vccd1 _18731_/Q sky130_fd_sc_hd__dfxtp_1
X_11066_ _10807_/A _11063_/X _11065_/X _10793_/A vssd1 vssd1 vccd1 vccd1 _11066_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15943_ _15943_/A vssd1 vssd1 vccd1 vccd1 _18972_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10017_ _10020_/A _10014_/X _10016_/X _09988_/X vssd1 vssd1 vccd1 vccd1 _10017_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18662_ _19608_/CLK _18662_/D vssd1 vssd1 vccd1 vccd1 _18662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15874_ _15055_/X _18942_/Q _15874_/S vssd1 vssd1 vccd1 vccd1 _15875_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17613_ _17723_/A vssd1 vssd1 vccd1 vccd1 _17707_/A sky130_fd_sc_hd__clkbuf_2
X_14825_ _14825_/A vssd1 vssd1 vccd1 vccd1 _14838_/A sky130_fd_sc_hd__clkbuf_2
X_18593_ _18853_/CLK _18593_/D vssd1 vssd1 vccd1 vccd1 _18593_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12608__B2 _19677_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17544_ _19632_/Q _16755_/A _17546_/S vssd1 vssd1 vccd1 vccd1 _17545_/A sky130_fd_sc_hd__mux2_1
X_14756_ _14765_/A _14765_/C vssd1 vssd1 vccd1 vccd1 _14756_/X sky130_fd_sc_hd__xor2_1
X_11968_ _12480_/A _11967_/X _12005_/A vssd1 vssd1 vccd1 vccd1 _11969_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09312__A _10793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13707_ _13724_/B _13580_/B vssd1 vssd1 vccd1 vccd1 _13922_/A sky130_fd_sc_hd__or2b_2
XANTENNA__09580__S0 _09344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17475_ _17475_/A vssd1 vssd1 vccd1 vccd1 _19601_/D sky130_fd_sc_hd__clkbuf_1
X_10919_ _10959_/A vssd1 vssd1 vccd1 vccd1 _10919_/X sky130_fd_sc_hd__buf_4
X_14687_ _11517_/B _14633_/X _14680_/X input54/X vssd1 vssd1 vccd1 vccd1 _14688_/B
+ sky130_fd_sc_hd__a22o_1
X_11899_ _11899_/A _11899_/B vssd1 vssd1 vccd1 vccd1 _11899_/Y sky130_fd_sc_hd__xnor2_4
X_19214_ _19597_/CLK _19214_/D vssd1 vssd1 vccd1 vccd1 _19214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16426_ _19177_/Q _15586_/X _16428_/S vssd1 vssd1 vccd1 vccd1 _16427_/A sky130_fd_sc_hd__mux2_1
X_13638_ _13636_/X _13637_/X _13741_/S vssd1 vssd1 vccd1 vccd1 _13638_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19145_ _19713_/CLK _19145_/D vssd1 vssd1 vccd1 vccd1 _19145_/Q sky130_fd_sc_hd__dfxtp_1
X_16357_ _16919_/A _16357_/B _15412_/C vssd1 vssd1 vccd1 vccd1 _16992_/B sky130_fd_sc_hd__or3b_4
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13569_ _11474_/A _11471_/A _11474_/B _11599_/A _11599_/C vssd1 vssd1 vccd1 vccd1
+ _13573_/C sky130_fd_sc_hd__o311a_1
XFILLER_173_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14591__C input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15308_ _15308_/A vssd1 vssd1 vccd1 vccd1 _18706_/D sky130_fd_sc_hd__clkbuf_1
X_19076_ _19659_/CLK _19076_/D vssd1 vssd1 vccd1 vccd1 _19076_/Q sky130_fd_sc_hd__dfxtp_1
X_16288_ _16033_/X _19115_/Q _16296_/S vssd1 vssd1 vccd1 vccd1 _16289_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13336__A2 _13334_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18027_ _18027_/A _18031_/C vssd1 vssd1 vccd1 vccd1 _18027_/Y sky130_fd_sc_hd__nor2_1
XFILLER_161_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15239_ _18682_/Q _15238_/X _15239_/S vssd1 vssd1 vccd1 vccd1 _15240_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09982__A _10256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15195__S _15201_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09800_ _09217_/A _09788_/X _09790_/X _09799_/X _09249_/X vssd1 vssd1 vccd1 vccd1
+ _09800_/X sky130_fd_sc_hd__a311o_4
XFILLER_114_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_82_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19786_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12612__S _12628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09731_ _10132_/A _09727_/Y _09730_/Y _10182_/A vssd1 vssd1 vccd1 vccd1 _09731_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18929_ _19549_/CLK _18929_/D vssd1 vssd1 vccd1 vccd1 _18929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17235__A0 _18454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09662_ _09662_/A vssd1 vssd1 vccd1 vccd1 _10245_/A sky130_fd_sc_hd__buf_2
XFILLER_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_97_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19780_/CLK sky130_fd_sc_hd__clkbuf_16
X_09593_ _11186_/S vssd1 vssd1 vccd1 vccd1 _10185_/S sky130_fd_sc_hd__buf_4
XANTENNA__11752__A _19731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13272__A1 _19672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09222__A _19694_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19712_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10368__A _10368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__S1 _09610_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14221__B1 _15123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_35_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19551_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_136_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13398__B _13398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11199__A _11199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09892__A _09892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12838__A1 _12840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09929_ _09928_/A _09913_/Y _09928_/Y _09826_/A vssd1 vssd1 vccd1 vccd1 _09929_/Y
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__11646__B _12462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09703__A1 _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15833__S _15841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12940_ _12943_/A _12940_/B _12946_/C vssd1 vssd1 vccd1 vccd1 _18290_/D sky130_fd_sc_hd__nor3_1
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12871_ _12873_/B _12873_/C _12870_/Y vssd1 vssd1 vccd1 vccd1 _18270_/D sky130_fd_sc_hd__o21a_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ input60/X vssd1 vssd1 vccd1 vccd1 _14610_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11662__A _19730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15134__A _15134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _12545_/A _11822_/B _15263_/A _11822_/D vssd1 vssd1 vccd1 vccd1 _11822_/X
+ sky130_fd_sc_hd__or4_2
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _18816_/Q _15589_/X _15590_/S vssd1 vssd1 vccd1 vccd1 _15591_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10077__A1 _09173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09132__A _10373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11381__B _12555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11753_ _19731_/Q _11752_/C _19732_/Q vssd1 vssd1 vccd1 vccd1 _11754_/B sky130_fd_sc_hd__a21oi_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14541_ _16430_/A _14582_/B vssd1 vssd1 vccd1 vccd1 _14541_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10172__S1 _11189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10704_ _10694_/Y _10698_/Y _10701_/Y _10703_/Y _10944_/A vssd1 vssd1 vccd1 vccd1
+ _10705_/A sky130_fd_sc_hd__o221a_1
XFILLER_53_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _17317_/S vssd1 vssd1 vccd1 vccd1 _17269_/S sky130_fd_sc_hd__buf_2
X_11684_ _11684_/A _11684_/B vssd1 vssd1 vccd1 vccd1 _11685_/A sky130_fd_sc_hd__and2_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14472_ _18507_/Q _19745_/Q _14476_/S vssd1 vssd1 vccd1 vccd1 _14473_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16211_ _18207_/A _16211_/B vssd1 vssd1 vccd1 vccd1 _19082_/D sky130_fd_sc_hd__nor2_1
X_13423_ _12577_/X _13415_/Y _13422_/X _12596_/X _18649_/Q vssd1 vssd1 vccd1 vccd1
+ _13423_/X sky130_fd_sc_hd__a32o_4
X_10635_ _19605_/Q _19443_/Q _18889_/Q _18659_/Q _10631_/X _10634_/X vssd1 vssd1 vccd1
+ vccd1 _10636_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13589__A _14332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17191_ _18441_/Q _13307_/X _17201_/S vssd1 vssd1 vccd1 vccd1 _17191_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12774__B1 _12735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13354_ _13354_/A vssd1 vssd1 vccd1 vccd1 _13354_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16142_ _16033_/X _19046_/Q _16150_/S vssd1 vssd1 vccd1 vccd1 _16143_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10566_ _10566_/A _10566_/B vssd1 vssd1 vccd1 vccd1 _10566_/X sky130_fd_sc_hd__or2_1
XFILLER_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ _14265_/A _12305_/B vssd1 vssd1 vccd1 vccd1 _12310_/A sky130_fd_sc_hd__xor2_1
XANTENNA__13101__B _13104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13285_ _18281_/Q _13326_/B vssd1 vssd1 vccd1 vccd1 _13285_/X sky130_fd_sc_hd__and2_1
XFILLER_115_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16073_ _16073_/A vssd1 vssd1 vccd1 vccd1 _19025_/D sky130_fd_sc_hd__clkbuf_1
X_10497_ _19640_/Q _19057_/Q _19094_/Q _18700_/Q _10450_/S _10239_/A vssd1 vssd1 vccd1
+ vccd1 _10498_/B sky130_fd_sc_hd__mux4_2
XFILLER_142_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15024_ _15024_/A vssd1 vssd1 vccd1 vccd1 _18612_/D sky130_fd_sc_hd__clkbuf_1
X_12236_ _12181_/A _14203_/B _12210_/A vssd1 vssd1 vccd1 vccd1 _12237_/B sky130_fd_sc_hd__a21oi_1
XFILLER_142_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19832_ _19833_/CLK _19832_/D vssd1 vssd1 vccd1 vccd1 _19832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11837__A _13653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12167_ _11706_/X _12165_/X _12166_/X _12072_/X vssd1 vssd1 vccd1 vccd1 _12167_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11118_ _19514_/Q _19128_/Q _19578_/Q _18734_/Q _09583_/A _10390_/A vssd1 vssd1 vccd1
+ vccd1 _11119_/B sky130_fd_sc_hd__mux4_1
X_19763_ _19861_/CLK _19763_/D vssd1 vssd1 vccd1 vccd1 _19763_/Q sky130_fd_sc_hd__dfxtp_1
X_16975_ _16822_/X _19395_/Q _16975_/S vssd1 vssd1 vccd1 vccd1 _16976_/A sky130_fd_sc_hd__mux2_1
X_12098_ _19675_/Q _12098_/B vssd1 vssd1 vccd1 vccd1 _12098_/X sky130_fd_sc_hd__or2_1
XFILLER_1_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10460__B _12480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16839__S _16839_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18714_ _19721_/CLK _18714_/D vssd1 vssd1 vccd1 vccd1 _18714_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15743__S _15747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15926_ _15937_/A vssd1 vssd1 vccd1 vccd1 _15935_/S sky130_fd_sc_hd__buf_4
X_11049_ _11060_/A _11049_/B vssd1 vssd1 vccd1 vccd1 _11049_/X sky130_fd_sc_hd__or2_1
XFILLER_49_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19694_ _19695_/CLK _19694_/D vssd1 vssd1 vccd1 vccd1 _19694_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_83_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17768__A1 _12193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 io_dbus_rdata[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__10304__A2 _19098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18645_ _19727_/CLK _18645_/D vssd1 vssd1 vccd1 vccd1 _18645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15857_ _14964_/X _18934_/Q _15863_/S vssd1 vssd1 vccd1 vccd1 _15858_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14808_ _16771_/A vssd1 vssd1 vccd1 vccd1 _14808_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18576_ _18618_/CLK _18576_/D vssd1 vssd1 vccd1 vccd1 _18576_/Q sky130_fd_sc_hd__dfxtp_1
X_15788_ _15788_/A vssd1 vssd1 vccd1 vccd1 _18903_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12387__B _19756_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17527_ _19625_/Q _16731_/X _17529_/S vssd1 vssd1 vccd1 vccd1 _17528_/A sky130_fd_sc_hd__mux2_1
X_14739_ _16648_/A vssd1 vssd1 vccd1 vccd1 _16752_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11722__D _11822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17458_ _17458_/A vssd1 vssd1 vccd1 vccd1 _19594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16409_ _19169_/Q _15561_/X _16413_/S vssd1 vssd1 vccd1 vccd1 _16410_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17389_ _16844_/X _19564_/Q _17389_/S vssd1 vssd1 vccd1 vccd1 _17390_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19128_ _19546_/CLK _19128_/D vssd1 vssd1 vccd1 vccd1 _19128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14107__B _14111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15918__S _15924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19059_ _19546_/CLK _19059_/D vssd1 vssd1 vccd1 vccd1 _19059_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14822__S _14822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15219__A _16721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17208__A0 _18446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11179__S0 _09729_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09714_ _11168_/A _09714_/B vssd1 vssd1 vccd1 vccd1 _09714_/X sky130_fd_sc_hd__or2_1
XANTENNA__13493__A1 _13346_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10926__S0 _10668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09645_ _19270_/Q _19041_/Q _18972_/Q _19366_/Q _11153_/A _09636_/X vssd1 vssd1 vccd1
+ vccd1 _09645_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12578__A _12766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09576_ _10329_/A vssd1 vssd1 vccd1 vccd1 _10331_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13245__B2 _18628_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16484__S _16486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10420_ _09642_/A _10417_/X _10419_/X vssd1 vssd1 vccd1 vccd1 _10420_/X sky130_fd_sc_hd__a21o_1
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17695__A0 _19675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10351_ _09171_/A _10350_/X _10475_/A vssd1 vssd1 vccd1 vccd1 _10351_/X sky130_fd_sc_hd__a21o_1
XFILLER_164_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13070_ _18112_/D vssd1 vssd1 vccd1 vccd1 _18110_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10282_ _18769_/Q _18998_/Q _18929_/Q _19227_/Q _09342_/A _11113_/A vssd1 vssd1 vccd1
+ vccd1 _10282_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12021_ _11790_/A _12019_/Y _12075_/C _12116_/A vssd1 vssd1 vccd1 vccd1 _12021_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_3_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11731__A1 _19731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10090__S0 _10153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16659__S _16671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16760_ _16760_/A vssd1 vssd1 vccd1 vccd1 _19311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13484__A1 _12617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13972_ _13969_/S _13777_/X _13816_/A vssd1 vssd1 vccd1 vccd1 _13972_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_76_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15711_ _18869_/Q _15554_/X _15719_/S vssd1 vssd1 vccd1 vccd1 _15712_/A sky130_fd_sc_hd__mux2_1
X_12923_ _12930_/C _12930_/D _12922_/X vssd1 vssd1 vccd1 vccd1 _12923_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16691_ _19290_/Q _16689_/X _16703_/S vssd1 vssd1 vccd1 vccd1 _16692_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12488__A _12488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10393__S1 _11111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18430_ _19691_/CLK _18430_/D vssd1 vssd1 vccd1 vccd1 _18430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15642_ _15642_/A vssd1 vssd1 vccd1 vccd1 _18838_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _18266_/Q _18265_/Q _18264_/Q _12854_/D vssd1 vssd1 vccd1 vccd1 _12865_/D
+ sky130_fd_sc_hd__and4_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _19082_/CLK _18361_/D vssd1 vssd1 vccd1 vccd1 _18361_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _12468_/A _12005_/A _11911_/C _14578_/A vssd1 vssd1 vccd1 vccd1 _13984_/A
+ sky130_fd_sc_hd__a2bb2o_4
X_15573_ _15573_/A vssd1 vssd1 vccd1 vccd1 _18810_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output100_A _11787_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16394__S _16402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18175__A _19845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12785_ _16212_/A _16138_/B vssd1 vssd1 vccd1 vccd1 _15413_/A sky130_fd_sc_hd__or2_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10145__S1 _09595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _17312_/A vssd1 vssd1 vccd1 vccd1 _19529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14524_ _14524_/A _14551_/B vssd1 vssd1 vccd1 vccd1 _14524_/Y sky130_fd_sc_hd__nand2_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18292_ _18298_/CLK _18292_/D vssd1 vssd1 vccd1 vccd1 _18292_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11736_ _11736_/A _11736_/B _11736_/C vssd1 vssd1 vccd1 vccd1 _11736_/X sky130_fd_sc_hd__or3_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17243_ _17243_/A vssd1 vssd1 vccd1 vccd1 _19499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14455_ _14455_/A vssd1 vssd1 vccd1 vccd1 _18499_/D sky130_fd_sc_hd__clkbuf_1
X_11667_ _12411_/B _11667_/B vssd1 vssd1 vccd1 vccd1 _11667_/X sky130_fd_sc_hd__and2b_1
XANTENNA__13112__A _13112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12654__C _14946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13406_ _19688_/Q _12737_/A _13205_/A _18412_/Q vssd1 vssd1 vccd1 vccd1 _13407_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17174_ _18436_/Q _13259_/X _17184_/S vssd1 vssd1 vccd1 vccd1 _17174_/X sky130_fd_sc_hd__mux2_1
X_10618_ _10873_/A _10618_/B vssd1 vssd1 vccd1 vccd1 _10618_/X sky130_fd_sc_hd__or2_1
X_11598_ _11639_/A _11598_/B vssd1 vssd1 vccd1 vccd1 _11686_/A sky130_fd_sc_hd__or2_1
X_14386_ _14386_/A vssd1 vssd1 vccd1 vccd1 _18473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17686__A0 _13307_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16125_ _16835_/A vssd1 vssd1 vccd1 vccd1 _16125_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13337_ _13390_/A _18641_/Q vssd1 vssd1 vccd1 vccd1 _13337_/Y sky130_fd_sc_hd__nand2_1
X_10549_ _18763_/Q _18992_/Q _18923_/Q _19221_/Q _10353_/A _10548_/X vssd1 vssd1 vccd1
+ vccd1 _10550_/B sky130_fd_sc_hd__mux4_1
XFILLER_128_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17150__A2 _17628_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16056_ _16055_/X _19020_/Q _16065_/S vssd1 vssd1 vccd1 vccd1 _16057_/A sky130_fd_sc_hd__mux2_1
X_13268_ _13324_/A vssd1 vssd1 vccd1 vccd1 _13403_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12670__B _14562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09915__A1 _09163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15007_ _14999_/X _15001_/X _15004_/Y _15006_/X vssd1 vssd1 vccd1 vccd1 _16721_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_155_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12219_ _14211_/A _12218_/X _12219_/S vssd1 vssd1 vccd1 vccd1 _12219_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13199_ _13438_/B vssd1 vssd1 vccd1 vccd1 _13246_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_124_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19815_ _19822_/CLK _19815_/D vssd1 vssd1 vccd1 vccd1 _19815_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10081__S0 _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14878__A _16686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16569__S _16569_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10930__C1 _09244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15473__S _15481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19746_ _19753_/CLK _19746_/D vssd1 vssd1 vccd1 vccd1 _19746_/Q sky130_fd_sc_hd__dfxtp_4
X_16958_ _16797_/X _19387_/Q _16964_/S vssd1 vssd1 vccd1 vccd1 _16959_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13475__A1 _13294_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15909_ _14856_/X _18957_/Q _15913_/S vssd1 vssd1 vccd1 vccd1 _15910_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19677_ _19680_/CLK _19677_/D vssd1 vssd1 vccd1 vccd1 _19677_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_65_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16889_ _19357_/Q _16699_/X _16891_/S vssd1 vssd1 vccd1 vccd1 _16890_/A sky130_fd_sc_hd__mux2_1
X_09430_ _09430_/A vssd1 vssd1 vccd1 vccd1 _09430_/X sky130_fd_sc_hd__buf_2
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18628_ _18632_/CLK _18628_/D vssd1 vssd1 vccd1 vccd1 _18628_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09361_ _09880_/A vssd1 vssd1 vccd1 vccd1 _09810_/A sky130_fd_sc_hd__buf_2
XFILLER_52_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09526__S0 _10242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18559_ _18585_/CLK _18559_/D vssd1 vssd1 vccd1 vccd1 _18559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18085__A _18085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_143_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09292_ _18531_/Q vssd1 vssd1 vccd1 vccd1 _15134_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14727__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14727__B2 _14711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17677__A0 _19672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12861__A _12991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput130 _12501_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[27] sky130_fd_sc_hd__buf_2
XFILLER_115_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput141 _12473_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[8] sky130_fd_sc_hd__buf_2
Xoutput152 _17888_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[17] sky130_fd_sc_hd__buf_2
XFILLER_115_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput163 _12370_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[27] sky130_fd_sc_hd__buf_2
Xoutput174 _17870_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[8] sky130_fd_sc_hd__buf_2
XFILLER_115_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_68_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09628_ _11200_/A _12503_/A vssd1 vssd1 vccd1 vccd1 _11220_/A sky130_fd_sc_hd__nand2_2
XFILLER_70_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09559_ _10417_/S vssd1 vssd1 vccd1 vccd1 _09700_/A sky130_fd_sc_hd__buf_2
XFILLER_102_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11940__A _11940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ _13440_/S vssd1 vssd1 vccd1 vccd1 _13092_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10452__A1 _10239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11521_ _11561_/A _13527_/C vssd1 vssd1 vccd1 vccd1 _11549_/A sky130_fd_sc_hd__and2_1
XFILLER_168_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11452_ _12715_/A _14718_/B vssd1 vssd1 vccd1 vccd1 _14431_/A sky130_fd_sc_hd__nand2_4
XANTENNA__13926__C1 _13711_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14240_ _14088_/X _14237_/Y _14239_/X vssd1 vssd1 vccd1 vccd1 _14240_/Y sky130_fd_sc_hd__o21ai_1
X_10403_ _10438_/A _10403_/B vssd1 vssd1 vccd1 vccd1 _10403_/Y sky130_fd_sc_hd__nor2_1
X_14171_ _14150_/X _14122_/X _14170_/X vssd1 vssd1 vccd1 vccd1 _14171_/X sky130_fd_sc_hd__a21o_1
XFILLER_164_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11383_ _11462_/A _13532_/A vssd1 vssd1 vccd1 vccd1 _12715_/A sky130_fd_sc_hd__nor2_2
XFILLER_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input61_A io_ibus_inst[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ _13171_/A _18619_/Q vssd1 vssd1 vccd1 vccd1 _13122_/Y sky130_fd_sc_hd__nand2_1
X_10334_ _10325_/A _10329_/X _10331_/Y _10333_/Y vssd1 vssd1 vccd1 vccd1 _10334_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_124_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17930_ _19761_/Q _17926_/C _17929_/Y vssd1 vssd1 vccd1 vccd1 _19761_/D sky130_fd_sc_hd__o21a_1
XFILLER_152_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13053_ _13055_/A _13055_/C _13052_/Y vssd1 vssd1 vccd1 vccd1 _18328_/D sky130_fd_sc_hd__o21a_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10265_ _19517_/Q _19131_/Q _19581_/Q _18737_/Q _09794_/A _09697_/A vssd1 vssd1 vccd1
+ vccd1 _10266_/B sky130_fd_sc_hd__mux4_1
XFILLER_133_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12004_ _11941_/Y _11282_/A _12026_/A vssd1 vssd1 vccd1 vccd1 _12004_/X sky130_fd_sc_hd__mux2_1
X_17861_ _17861_/A vssd1 vssd1 vccd1 vccd1 _19731_/D sky130_fd_sc_hd__clkbuf_1
X_10196_ _10196_/A _12487_/A vssd1 vssd1 vccd1 vccd1 _10197_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14698__A _17890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16389__S _16391_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16812_ _16812_/A vssd1 vssd1 vccd1 vccd1 _19327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16643__A1 _16639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19600_ _19699_/CLK _19600_/D vssd1 vssd1 vccd1 vccd1 _19600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17792_ _15149_/X _19699_/Q _17794_/S vssd1 vssd1 vccd1 vccd1 _17793_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19531_ _19713_/CLK _19531_/D vssd1 vssd1 vccd1 vccd1 _19531_/Q sky130_fd_sc_hd__dfxtp_1
X_16743_ _16743_/A vssd1 vssd1 vccd1 vccd1 _16743_/X sky130_fd_sc_hd__buf_2
X_13955_ _13993_/A _13955_/B vssd1 vssd1 vccd1 vccd1 _13955_/X sky130_fd_sc_hd__or2_1
XFILLER_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12906_ _17999_/A vssd1 vssd1 vccd1 vccd1 _12997_/A sky130_fd_sc_hd__buf_4
XFILLER_35_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19462_ _19592_/CLK _19462_/D vssd1 vssd1 vccd1 vccd1 _19462_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13209__A1 _19830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12011__A _12011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16674_ _16741_/S vssd1 vssd1 vccd1 vccd1 _16687_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_34_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09304__B _09624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13886_ _13884_/X _13885_/X _13965_/S vssd1 vssd1 vccd1 vccd1 _13886_/X sky130_fd_sc_hd__mux2_1
X_18413_ _19791_/CLK _18413_/D vssd1 vssd1 vccd1 vccd1 _18413_/Q sky130_fd_sc_hd__dfxtp_1
X_15625_ _18831_/Q _15535_/X _15625_/S vssd1 vssd1 vccd1 vccd1 _15626_/A sky130_fd_sc_hd__mux2_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _12840_/B _12840_/C _12817_/X vssd1 vssd1 vccd1 vccd1 _12837_/Y sky130_fd_sc_hd__a21oi_1
X_19393_ _19587_/CLK _19393_/D vssd1 vssd1 vccd1 vccd1 _19393_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10691__B2 _18433_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12946__A _18292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _19759_/CLK _18344_/D vssd1 vssd1 vccd1 vccd1 _18344_/Q sky130_fd_sc_hd__dfxtp_1
X_15556_ _18805_/Q _15554_/X _15568_/S vssd1 vssd1 vccd1 vccd1 _15557_/A sky130_fd_sc_hd__mux2_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _13154_/B vssd1 vssd1 vccd1 vccd1 _12768_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16137__B _16357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _14507_/A vssd1 vssd1 vccd1 vccd1 _18522_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18275_ _18386_/CLK _18275_/D vssd1 vssd1 vccd1 vccd1 _18275_/Q sky130_fd_sc_hd__dfxtp_1
X_11719_ _13166_/A _11719_/B vssd1 vssd1 vccd1 vccd1 _11726_/A sky130_fd_sc_hd__nand2_1
X_15487_ _16743_/A vssd1 vssd1 vccd1 vccd1 _15487_/X sky130_fd_sc_hd__buf_2
X_12699_ _14648_/A vssd1 vssd1 vccd1 vccd1 _13106_/B sky130_fd_sc_hd__buf_4
XFILLER_174_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17226_ _17226_/A vssd1 vssd1 vccd1 vccd1 _17239_/S sky130_fd_sc_hd__buf_2
Xinput10 io_dbus_rdata[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_4
X_14438_ _14438_/A vssd1 vssd1 vccd1 vccd1 _18491_/D sky130_fd_sc_hd__clkbuf_1
Xinput21 io_dbus_rdata[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_2
Xinput32 io_dbus_rdata[9] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__buf_2
XFILLER_156_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput43 io_ibus_inst[18] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_2
Xinput54 io_ibus_inst[28] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__buf_2
XANTENNA__15468__S _15470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17157_ _18431_/Q _13197_/X _17167_/S vssd1 vssd1 vccd1 vccd1 _17157_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14590__C1 _14585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17249__A _17317_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput65 io_ibus_inst[9] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_1
X_14369_ _14384_/A vssd1 vssd1 vccd1 vccd1 _14381_/S sky130_fd_sc_hd__clkbuf_2
X_16108_ _16108_/A vssd1 vssd1 vccd1 vccd1 _19036_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17088_ _17134_/S vssd1 vssd1 vccd1 vccd1 _17097_/S sky130_fd_sc_hd__buf_4
XFILLER_170_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16039_ _16749_/A vssd1 vssd1 vccd1 vccd1 _16039_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19729_ _19738_/CLK _19729_/D vssd1 vssd1 vccd1 vccd1 _19729_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__11744__B _11784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12120__A1 _19676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15931__S _15935_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10252__A1_N _18443_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ _09616_/A vssd1 vssd1 vccd1 vccd1 _09414_/A sky130_fd_sc_hd__buf_2
XFILLER_41_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14948__A1 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15070__B1 _14893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10109__S1 _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15232__A _16734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ _09344_/A vssd1 vssd1 vccd1 vccd1 _10055_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09230__A _09230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09275_ _09275_/A vssd1 vssd1 vccd1 vccd1 _09276_/A sky130_fd_sc_hd__buf_2
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15373__A1 _15184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15378__S _15384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10293__S0 _09675_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17593__S _17601_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10315__S _11157_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11000__A _18427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10045__S0 _09866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ _09927_/X _10040_/X _10049_/X _09309_/X _18447_/Q vssd1 vssd1 vccd1 vccd1
+ _12491_/C sky130_fd_sc_hd__a32o_4
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09738__S0 _09729_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15841__S _15841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13740_ _13997_/S vssd1 vssd1 vccd1 vccd1 _13913_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10122__B1 _09988_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ _10946_/A _10951_/X _10728_/X vssd1 vssd1 vccd1 vccd1 _10952_/X sky130_fd_sc_hd__o21a_1
XFILLER_90_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13671_ _13671_/A vssd1 vssd1 vccd1 vccd1 _13800_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10673__B2 _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12766__A _12766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10883_ _10895_/A _10883_/B vssd1 vssd1 vccd1 vccd1 _10883_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11670__A _19661_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15410_ _18752_/Q _15238_/X _15410_/S vssd1 vssd1 vccd1 vccd1 _15411_/A sky130_fd_sc_hd__mux2_1
X_12622_ _14562_/A _12622_/B vssd1 vssd1 vccd1 vccd1 _13236_/A sky130_fd_sc_hd__nor2_4
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16390_ _16390_/A vssd1 vssd1 vccd1 vccd1 _19160_/D sky130_fd_sc_hd__clkbuf_1
X_15341_ _15397_/A vssd1 vssd1 vccd1 vccd1 _15410_/S sky130_fd_sc_hd__buf_8
X_12553_ _18067_/B _12518_/X _12522_/X _13024_/B _12552_/X vssd1 vssd1 vccd1 vccd1
+ _12554_/B sky130_fd_sc_hd__a221o_2
XFILLER_106_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18060_ _18059_/A _18059_/C _19806_/Q vssd1 vssd1 vccd1 vccd1 _18061_/C sky130_fd_sc_hd__a21oi_1
X_11504_ _11519_/A _11519_/B _11519_/D vssd1 vssd1 vccd1 vccd1 _11512_/A sky130_fd_sc_hd__or3_1
XFILLER_11_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15272_ _18690_/Q _15143_/X _15278_/S vssd1 vssd1 vccd1 vccd1 _15273_/A sky130_fd_sc_hd__mux2_1
X_12484_ _12505_/B vssd1 vssd1 vccd1 vccd1 _12497_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_156_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17011_ _17011_/A vssd1 vssd1 vccd1 vccd1 _19410_/D sky130_fd_sc_hd__clkbuf_1
X_14223_ _14227_/A _14227_/B vssd1 vssd1 vccd1 vccd1 _14223_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11435_ _18419_/Q _12555_/B _18417_/Q vssd1 vssd1 vccd1 vccd1 _12557_/A sky130_fd_sc_hd__nor3b_2
XFILLER_7_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14154_ _13927_/X _14151_/Y _14153_/X _14003_/X vssd1 vssd1 vccd1 vccd1 _14154_/X
+ sky130_fd_sc_hd__a211o_1
X_11366_ _11366_/A _11366_/B _13584_/C _11365_/X vssd1 vssd1 vccd1 vccd1 _11367_/D
+ sky130_fd_sc_hd__or4b_1
XFILLER_153_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13105_ _18346_/Q _12731_/A _13104_/X _13102_/X vssd1 vssd1 vccd1 vccd1 _18346_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10317_ _10080_/X _10314_/X _10316_/X vssd1 vssd1 vccd1 vccd1 _10317_/X sky130_fd_sc_hd__a21o_1
X_11297_ _14511_/A _11297_/B _11297_/C vssd1 vssd1 vccd1 vccd1 _11298_/B sky130_fd_sc_hd__and3_1
XANTENNA__13678__A1 _14057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14085_ _13914_/X _13916_/X _14085_/S vssd1 vssd1 vccd1 vccd1 _14085_/X sky130_fd_sc_hd__mux2_1
X_18962_ _19645_/CLK _18962_/D vssd1 vssd1 vccd1 vccd1 _18962_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10036__S0 _09866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13036_ _13047_/D vssd1 vssd1 vccd1 vccd1 _13045_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_140_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17913_ _19792_/Q _19793_/Q _19795_/Q _19794_/Q vssd1 vssd1 vccd1 vccd1 _18026_/A
+ sky130_fd_sc_hd__and4_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ _10395_/A _10247_/X _09681_/A vssd1 vssd1 vccd1 vccd1 _10248_/X sky130_fd_sc_hd__o21a_1
X_18893_ _19223_/CLK _18893_/D vssd1 vssd1 vccd1 vccd1 _18893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17008__S _17014_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14859__C _14859_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17844_ _17844_/A vssd1 vssd1 vccd1 vccd1 _19722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10179_ _10175_/A _10178_/X _09616_/X vssd1 vssd1 vccd1 vccd1 _10179_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_113_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09315__A _09315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17775_ _17779_/A _17775_/B vssd1 vssd1 vccd1 vccd1 _17776_/A sky130_fd_sc_hd__and2_2
X_14987_ _14986_/X _18609_/Q _14997_/S vssd1 vssd1 vccd1 vccd1 _14988_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12102__A1 _17711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16726_ _19301_/Q _16725_/X _16735_/S vssd1 vssd1 vccd1 vccd1 _16727_/A sky130_fd_sc_hd__mux2_1
X_19514_ _19709_/CLK _19514_/D vssd1 vssd1 vccd1 vccd1 _19514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13938_ _14274_/A vssd1 vssd1 vccd1 vccd1 _14178_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19445_ _19639_/CLK _19445_/D vssd1 vssd1 vccd1 vccd1 _19445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16657_ _16657_/A vssd1 vssd1 vccd1 vccd1 _16657_/X sky130_fd_sc_hd__clkbuf_2
X_13869_ _13821_/A _13855_/Y _13868_/Y _13738_/X vssd1 vssd1 vccd1 vccd1 _13869_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15052__B1 _14842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15608_ _18823_/Q _15510_/X _15614_/S vssd1 vssd1 vccd1 vccd1 _15609_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19376_ _19569_/CLK _19376_/D vssd1 vssd1 vccd1 vccd1 _19376_/Q sky130_fd_sc_hd__dfxtp_1
X_16588_ _16588_/A vssd1 vssd1 vccd1 vccd1 _19249_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_16_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18327_ _19822_/CLK _18327_/D vssd1 vssd1 vccd1 vccd1 _18327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15539_ _15571_/A vssd1 vssd1 vccd1 vccd1 _15552_/S sky130_fd_sc_hd__buf_4
XANTENNA__10196__A _10196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18258_ _19855_/CLK _18258_/D vssd1 vssd1 vccd1 vccd1 _18258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17209_ _17226_/A vssd1 vssd1 vccd1 vccd1 _17223_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__15198__S _15201_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18189_ _19850_/Q _18191_/C _18188_/Y vssd1 vssd1 vccd1 vccd1 _19850_/D sky130_fd_sc_hd__o21a_1
XFILLER_144_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11916__A1 _18500_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10275__S0 _09675_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15107__A1 _18631_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15107__B2 _10461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09990__C1 _09854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09962_ _09385_/A _09961_/X _09319_/A vssd1 vssd1 vccd1 vccd1 _09962_/X sky130_fd_sc_hd__o21a_1
XFILLER_131_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09968__S0 _09872_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09893_ _09944_/A _09891_/X _09892_/X vssd1 vssd1 vccd1 vccd1 _09893_/Y sky130_fd_sc_hd__o21ai_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11852__A0 _11846_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16791__A0 _16790_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17588__S _17590_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09327_ _10496_/A vssd1 vssd1 vccd1 vccd1 _10288_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_138_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09258_ _18532_/Q vssd1 vssd1 vccd1 vccd1 _14716_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_138_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09189_ _10115_/A _09174_/X _09237_/A vssd1 vssd1 vccd1 vccd1 _09189_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11220_ _11220_/A _11220_/B vssd1 vssd1 vccd1 vccd1 _11220_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10040__C1 _09404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11151_ _11151_/A _11225_/A _11151_/C vssd1 vssd1 vccd1 vccd1 _11152_/D sky130_fd_sc_hd__and3_1
XFILLER_161_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10102_ _10102_/A _10102_/B vssd1 vssd1 vccd1 vccd1 _11227_/A sky130_fd_sc_hd__nor2_1
XFILLER_122_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09959__S0 _09872_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14321__A2 _14324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11082_ _12478_/B _11082_/B vssd1 vssd1 vccd1 vccd1 _11083_/A sky130_fd_sc_hd__and2b_1
XFILLER_103_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10033_ _18607_/Q _19296_/Q _10033_/S vssd1 vssd1 vccd1 vccd1 _10033_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10569__S1 _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14910_ _14910_/A vssd1 vssd1 vccd1 vccd1 _18602_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11665__A _19730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15137__A _16503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15890_ _15890_/A vssd1 vssd1 vccd1 vccd1 _18948_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10343__B1 _09317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09135__A _09135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A io_dbus_rdata[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14841_ _17662_/A _14840_/B _14829_/B vssd1 vssd1 vccd1 vccd1 _14841_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_124_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17560_ _19639_/Q _16777_/A _17568_/S vssd1 vssd1 vccd1 vccd1 _17561_/A sky130_fd_sc_hd__mux2_1
X_14772_ _16761_/A vssd1 vssd1 vccd1 vccd1 _14772_/X sky130_fd_sc_hd__buf_2
XFILLER_91_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11984_ _11984_/A _19739_/Q _17878_/A _11984_/D vssd1 vssd1 vccd1 vccd1 _12067_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_17_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16511_ _16511_/A vssd1 vssd1 vccd1 vccd1 _19213_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18220__B1 _12948_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13723_ _12511_/A _13806_/A _13711_/Y _13722_/X vssd1 vssd1 vccd1 vccd1 _13723_/X
+ sky130_fd_sc_hd__o211a_1
X_17491_ _17491_/A vssd1 vssd1 vccd1 vccd1 _19608_/D sky130_fd_sc_hd__clkbuf_1
X_10935_ _10772_/X _10934_/X _11062_/A vssd1 vssd1 vccd1 vccd1 _10935_/X sky130_fd_sc_hd__a21o_1
XFILLER_16_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19230_ _19326_/CLK _19230_/D vssd1 vssd1 vccd1 vccd1 _19230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16442_ _16048_/X _19183_/Q _16442_/S vssd1 vssd1 vccd1 vccd1 _16443_/A sky130_fd_sc_hd__mux2_1
X_13654_ _14034_/S vssd1 vssd1 vccd1 vccd1 _13995_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_32_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10866_ _10866_/A _10866_/B vssd1 vssd1 vccd1 vccd1 _10866_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ _18285_/Q vssd1 vssd1 vccd1 vccd1 _12930_/C sky130_fd_sc_hd__clkbuf_2
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19161_ _19223_/CLK _19161_/D vssd1 vssd1 vccd1 vccd1 _19161_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13104__B _13104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16373_ _16373_/A vssd1 vssd1 vccd1 vccd1 _19152_/D sky130_fd_sc_hd__clkbuf_1
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13585_ _13585_/A _13585_/B _13585_/C _13585_/D vssd1 vssd1 vccd1 vccd1 _13585_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__18183__A _19848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10797_ _10797_/A _10797_/B vssd1 vssd1 vccd1 vccd1 _10797_/X sky130_fd_sc_hd__or2_1
X_18112_ _19825_/Q _19824_/Q _18334_/Q _18112_/D vssd1 vssd1 vccd1 vccd1 _18122_/D
+ sky130_fd_sc_hd__and4_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15324_ _15324_/A vssd1 vssd1 vccd1 vccd1 _15333_/S sky130_fd_sc_hd__buf_4
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12536_ _12587_/A vssd1 vssd1 vccd1 vccd1 _12742_/A sky130_fd_sc_hd__buf_2
XFILLER_118_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19092_ _19638_/CLK _19092_/D vssd1 vssd1 vccd1 vccd1 _19092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18043_ _18043_/A _19800_/Q _18043_/C vssd1 vssd1 vccd1 vccd1 _18045_/B sky130_fd_sc_hd__and3_1
XFILLER_172_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15255_ _15255_/A _15255_/B vssd1 vssd1 vccd1 vccd1 _15255_/X sky130_fd_sc_hd__or2_1
XFILLER_145_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12467_ _12467_/A vssd1 vssd1 vccd1 vccd1 _12467_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__14216__A _14216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14206_ _13971_/X _14072_/X _14205_/X vssd1 vssd1 vccd1 vccd1 _14206_/X sky130_fd_sc_hd__a21o_1
X_11418_ _12520_/A _12751_/D _11419_/C vssd1 vssd1 vccd1 vccd1 _12585_/A sky130_fd_sc_hd__nor3_2
XFILLER_144_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15186_ _15186_/A vssd1 vssd1 vccd1 vccd1 _18665_/D sky130_fd_sc_hd__clkbuf_1
X_12398_ _13712_/A _14300_/A _12379_/B vssd1 vssd1 vccd1 vccd1 _12399_/B sky130_fd_sc_hd__a21bo_1
XFILLER_98_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09972__C1 _09395_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14137_ _13810_/X _13706_/B _14136_/X vssd1 vssd1 vccd1 vccd1 _14137_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_141_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11349_ _18585_/Q _11361_/A _11358_/B _13526_/C vssd1 vssd1 vccd1 vccd1 _11598_/B
+ sky130_fd_sc_hd__or4_2
XANTENNA__16431__A _16920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18945_ _19632_/CLK _18945_/D vssd1 vssd1 vccd1 vccd1 _18945_/Q sky130_fd_sc_hd__dfxtp_1
X_14068_ _11926_/Y _13827_/X _14067_/X _13828_/X vssd1 vssd1 vccd1 vccd1 _14068_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_86_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13019_ _13049_/A _13024_/C vssd1 vssd1 vccd1 vccd1 _13019_/Y sky130_fd_sc_hd__nor2_1
X_18876_ _19643_/CLK _18876_/D vssd1 vssd1 vccd1 vccd1 _18876_/Q sky130_fd_sc_hd__dfxtp_1
X_17827_ _15200_/X _19715_/Q _17827_/S vssd1 vssd1 vccd1 vccd1 _17828_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15481__S _15481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12626__A2 _12703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17758_ _17765_/C _17757_/Y _17713_/X vssd1 vssd1 vccd1 vccd1 _17758_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_82_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16709_ _16709_/A vssd1 vssd1 vccd1 vccd1 _16709_/X sky130_fd_sc_hd__clkbuf_2
X_17689_ _17689_/A vssd1 vssd1 vccd1 vccd1 _19674_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19428_ _19556_/CLK _19428_/D vssd1 vssd1 vccd1 vccd1 _19428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19359_ _19810_/CLK _19359_/D vssd1 vssd1 vccd1 vccd1 _19359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09112_ _11472_/A _11365_/B vssd1 vssd1 vccd1 vccd1 _09113_/B sky130_fd_sc_hd__nand2_4
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14126__A _14126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_13_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_116_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15656__S _15658_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09963__C1 _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14839__A0 _18437_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09945_ _18840_/Q _19394_/Q _19556_/Q _18808_/Q _09809_/X _09881_/X vssd1 vssd1 vccd1
+ vccd1 _09945_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09876_ _09826_/A _09873_/Y _09875_/Y _09947_/A vssd1 vssd1 vccd1 vccd1 _09876_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_112_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15391__S _15395_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12078__B1 _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10720_ _18760_/Q _18989_/Q _18920_/Q _19218_/Q _10719_/X _09481_/A vssd1 vssd1 vccd1
+ vccd1 _10721_/B sky130_fd_sc_hd__mux4_2
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_191_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _10651_/A _10651_/B vssd1 vssd1 vccd1 vccd1 _10651_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16516__A _16573_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17111__S _17119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11053__A1 _10713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13370_ _19685_/Q _12737_/X _15242_/D _18409_/Q vssd1 vssd1 vccd1 vccd1 _13370_/X
+ sky130_fd_sc_hd__a22o_1
X_10582_ _10238_/A _10581_/X _10638_/A vssd1 vssd1 vccd1 vccd1 _10582_/X sky130_fd_sc_hd__a21o_1
XFILLER_70_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12321_ _17711_/A _12319_/Y _12341_/B _17886_/A vssd1 vssd1 vccd1 vccd1 _12321_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_103_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15040_ _18454_/Q _13398_/B _15051_/S vssd1 vssd1 vccd1 vccd1 _15040_/X sky130_fd_sc_hd__mux2_1
X_12252_ _11790_/A _12250_/Y _12251_/X _12116_/A vssd1 vssd1 vccd1 vccd1 _12252_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_135_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11203_ _11203_/A _11203_/B vssd1 vssd1 vccd1 vccd1 _11249_/A sky130_fd_sc_hd__or2_2
X_12183_ _12138_/A _12161_/A _12161_/B vssd1 vssd1 vccd1 vccd1 _12183_/X sky130_fd_sc_hd__o21ba_1
XFILLER_122_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11134_ _11242_/A _11242_/B _11242_/C _11132_/Y _11133_/Y vssd1 vssd1 vccd1 vccd1
+ _11262_/B sky130_fd_sc_hd__a41o_1
XFILLER_96_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16991_ _16991_/A vssd1 vssd1 vccd1 vccd1 _19402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11065_ _11065_/A _11065_/B vssd1 vssd1 vccd1 vccd1 _11065_/X sky130_fd_sc_hd__or2_1
X_18730_ _19659_/CLK _18730_/D vssd1 vssd1 vccd1 vccd1 _18730_/Q sky130_fd_sc_hd__dfxtp_1
X_15942_ _15033_/X _18972_/Q _15946_/S vssd1 vssd1 vccd1 vccd1 _15943_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10316__B1 _09184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17244__A1 _18457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ _10074_/A _10016_/B vssd1 vssd1 vccd1 vccd1 _10016_/X sky130_fd_sc_hd__or2_1
XFILLER_76_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18661_ _19543_/CLK _18661_/D vssd1 vssd1 vccd1 vccd1 _18661_/Q sky130_fd_sc_hd__dfxtp_1
X_15873_ _15873_/A vssd1 vssd1 vccd1 vccd1 _18941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17612_ _12737_/X _15241_/X _17611_/Y _15243_/Y vssd1 vssd1 vccd1 vccd1 _17723_/A
+ sky130_fd_sc_hd__o211a_1
X_14824_ _14873_/A _14824_/B _14824_/C _14824_/D vssd1 vssd1 vccd1 vccd1 _14824_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_48_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18592_ _19704_/CLK _18592_/D vssd1 vssd1 vccd1 vccd1 _18592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11816__A0 _11813_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17543_ _17543_/A vssd1 vssd1 vccd1 vccd1 _19631_/D sky130_fd_sc_hd__clkbuf_1
X_14755_ _14755_/A vssd1 vssd1 vccd1 vccd1 _18589_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11842__B _13658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11967_ _11941_/Y _14543_/A _12026_/A vssd1 vssd1 vccd1 vccd1 _11967_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10739__A _10739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13706_ _13706_/A _13706_/B vssd1 vssd1 vccd1 vccd1 _13706_/Y sky130_fd_sc_hd__nor2_1
X_17474_ _19601_/Q _16654_/X _17474_/S vssd1 vssd1 vccd1 vccd1 _17475_/A sky130_fd_sc_hd__mux2_1
X_10918_ _19693_/Q vssd1 vssd1 vccd1 vccd1 _11026_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_1_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19708_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09580__S1 _11189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14686_ _14686_/A vssd1 vssd1 vccd1 vccd1 _18581_/D sky130_fd_sc_hd__clkbuf_1
X_11898_ _11879_/A _11879_/B _11871_/A vssd1 vssd1 vccd1 vccd1 _11899_/B sky130_fd_sc_hd__a21boi_2
XFILLER_20_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19213_ _19698_/CLK _19213_/D vssd1 vssd1 vccd1 vccd1 _19213_/Q sky130_fd_sc_hd__dfxtp_1
X_16425_ _16425_/A vssd1 vssd1 vccd1 vccd1 _19176_/D sky130_fd_sc_hd__clkbuf_1
X_13637_ _11843_/A _12307_/A _13657_/S vssd1 vssd1 vccd1 vccd1 _13637_/X sky130_fd_sc_hd__mux2_1
X_10849_ _19506_/Q _19120_/Q _19570_/Q _18726_/Q _10648_/S _10634_/A vssd1 vssd1 vccd1
+ vccd1 _10850_/B sky130_fd_sc_hd__mux4_1
XFILLER_60_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17021__S _17025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19144_ _19725_/CLK _19144_/D vssd1 vssd1 vccd1 vccd1 _19144_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10478__S0 _09447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16356_ _16356_/A vssd1 vssd1 vccd1 vccd1 _19146_/D sky130_fd_sc_hd__clkbuf_1
X_13568_ _13568_/A _13568_/B vssd1 vssd1 vccd1 vccd1 _13573_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15307_ _18706_/Q _15194_/X _15311_/S vssd1 vssd1 vccd1 vccd1 _15308_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12519_ _12519_/A vssd1 vssd1 vccd1 vccd1 _12791_/A sky130_fd_sc_hd__buf_2
X_19075_ _19724_/CLK _19075_/D vssd1 vssd1 vccd1 vccd1 _19075_/Q sky130_fd_sc_hd__dfxtp_1
X_16287_ _16355_/S vssd1 vssd1 vccd1 vccd1 _16296_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_173_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13499_ _13499_/A vssd1 vssd1 vccd1 vccd1 _13508_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18026_ _18026_/A vssd1 vssd1 vccd1 vccd1 _18031_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15238_ _16740_/A vssd1 vssd1 vccd1 vccd1 _15238_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15169_ _18660_/Q _15168_/X _15169_/S vssd1 vssd1 vccd1 vccd1 _15170_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09730_ _09867_/A _09730_/B vssd1 vssd1 vccd1 vccd1 _09730_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18928_ _19549_/CLK _18928_/D vssd1 vssd1 vccd1 vccd1 _18928_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10307__A0 _19612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17235__A1 _13399_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10402__S0 _11112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09661_ _09661_/A _09661_/B vssd1 vssd1 vccd1 vccd1 _09661_/Y sky130_fd_sc_hd__nor2_1
X_18859_ _19543_/CLK _18859_/D vssd1 vssd1 vccd1 vccd1 _18859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09592_ _09675_/S vssd1 vssd1 vccd1 vccd1 _11186_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_39_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11752__B _19732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11807__B1 _11970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13025__A _13034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12864__A _12904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11035__A1 _10821_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10469__S0 _09447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17171__A0 _18435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10384__A _10384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11199__B _12502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10641__S0 _10631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_138_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12299__B1 _17241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09928_ _09928_/A _18872_/Q vssd1 vssd1 vccd1 vccd1 _09928_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09859_ _18842_/Q _19396_/Q _19558_/Q _18810_/Q _09163_/A _09843_/A vssd1 vssd1 vccd1
+ vccd1 _09859_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17106__S _17108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15415__A _16503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12870_ _12873_/B _12873_/C _12869_/X vssd1 vssd1 vccd1 vccd1 _12870_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16010__S _16016_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _11821_/A vssd1 vssd1 vccd1 vccd1 _12545_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11662__B _13529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16945__S _16953_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10559__A _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _15339_/A vssd1 vssd1 vccd1 vccd1 _16430_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_14_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11752_ _19731_/Q _19732_/Q _11752_/C vssd1 vssd1 vccd1 vccd1 _11792_/B sky130_fd_sc_hd__and3_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10482__C1 _09246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10703_ _10791_/A _10702_/X _10793_/A vssd1 vssd1 vccd1 vccd1 _10703_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _14471_/A vssd1 vssd1 vccd1 vccd1 _18506_/D sky130_fd_sc_hd__clkbuf_1
X_11683_ _17143_/S _11668_/X _11670_/X _11682_/Y _11997_/A vssd1 vssd1 vccd1 vccd1
+ _11684_/B sky130_fd_sc_hd__a311o_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _16210_/A vssd1 vssd1 vccd1 vccd1 _19077_/D sky130_fd_sc_hd__clkbuf_1
X_13422_ _18649_/Q _13422_/B vssd1 vssd1 vccd1 vccd1 _13422_/X sky130_fd_sc_hd__or2_1
X_17190_ _17190_/A vssd1 vssd1 vccd1 vccd1 _19483_/D sky130_fd_sc_hd__clkbuf_1
X_10634_ _10634_/A vssd1 vssd1 vccd1 vccd1 _10634_/X sky130_fd_sc_hd__buf_4
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12493__B _12495_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16141_ _16209_/S vssd1 vssd1 vccd1 vccd1 _16150_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__12774__B2 _19848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13353_ _12779_/X _13139_/X _13352_/X _13350_/X vssd1 vssd1 vccd1 vccd1 _18374_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10565_ _18762_/Q _18991_/Q _18922_/Q _19220_/Q _10604_/S _10422_/A vssd1 vssd1 vccd1
+ vccd1 _10566_/B sky130_fd_sc_hd__mux4_1
XFILLER_5_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ _12256_/A _12258_/B _12280_/A _13567_/A vssd1 vssd1 vccd1 vccd1 _12305_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_115_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14515__A2 _12692_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16072_ _16071_/X _19025_/Q _16081_/S vssd1 vssd1 vccd1 vccd1 _16073_/A sky130_fd_sc_hd__mux2_1
X_13284_ _13403_/A _18633_/Q vssd1 vssd1 vccd1 vccd1 _13284_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10496_ _10496_/A _10496_/B vssd1 vssd1 vccd1 vccd1 _10496_/X sky130_fd_sc_hd__or2_1
XFILLER_154_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15023_ _15022_/X _18612_/Q _15056_/S vssd1 vssd1 vccd1 vccd1 _15024_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15296__S _15300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17077__A _17134_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12235_ _12235_/A vssd1 vssd1 vccd1 vccd1 _12235_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19831_ _19833_/CLK _19831_/D vssd1 vssd1 vccd1 vccd1 _19831_/Q sky130_fd_sc_hd__dfxtp_1
X_12166_ _19678_/Q _12390_/B vssd1 vssd1 vccd1 vccd1 _12166_/X sky130_fd_sc_hd__or2_1
XANTENNA__11837__B _13984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11117_ _10219_/X _11107_/Y _11109_/Y _09393_/A _11116_/X vssd1 vssd1 vccd1 vccd1
+ _11117_/X sky130_fd_sc_hd__o311a_2
X_19762_ _19861_/CLK _19762_/D vssd1 vssd1 vccd1 vccd1 _19762_/Q sky130_fd_sc_hd__dfxtp_1
X_16974_ _16974_/A vssd1 vssd1 vccd1 vccd1 _19394_/D sky130_fd_sc_hd__clkbuf_1
X_12097_ _12294_/S _12092_/X _12095_/Y _12096_/X _11980_/A vssd1 vssd1 vccd1 vccd1
+ _12097_/X sky130_fd_sc_hd__a311o_1
XFILLER_110_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18713_ _19718_/CLK _18713_/D vssd1 vssd1 vccd1 vccd1 _18713_/Q sky130_fd_sc_hd__dfxtp_1
X_15925_ _15925_/A vssd1 vssd1 vccd1 vccd1 _18964_/D sky130_fd_sc_hd__clkbuf_1
X_11048_ _19243_/Q _19014_/Q _18945_/Q _19339_/Q _10710_/A _10940_/X vssd1 vssd1 vccd1
+ vccd1 _11049_/B sky130_fd_sc_hd__mux4_2
XFILLER_83_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19693_ _19693_/CLK _19693_/D vssd1 vssd1 vccd1 vccd1 _19693_/Q sky130_fd_sc_hd__dfxtp_2
Xinput8 io_dbus_rdata[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XANTENNA__17768__A2 _13423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11853__A _19666_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15856_ _15856_/A vssd1 vssd1 vccd1 vccd1 _18933_/D sky130_fd_sc_hd__clkbuf_1
X_18644_ _19628_/CLK _18644_/D vssd1 vssd1 vccd1 vccd1 _18644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14807_ _16667_/A vssd1 vssd1 vccd1 vccd1 _16771_/A sky130_fd_sc_hd__clkbuf_2
X_15787_ _14975_/X _18903_/Q _15791_/S vssd1 vssd1 vccd1 vccd1 _15788_/A sky130_fd_sc_hd__mux2_1
X_18575_ _18618_/CLK _18575_/D vssd1 vssd1 vccd1 vccd1 _18575_/Q sky130_fd_sc_hd__dfxtp_2
X_12999_ _18313_/Q vssd1 vssd1 vccd1 vccd1 _13003_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14738_ _14732_/X _14736_/X _14737_/Y input23/X _14703_/X vssd1 vssd1 vccd1 vccd1
+ _16648_/A sky130_fd_sc_hd__a32o_1
X_17526_ _17526_/A vssd1 vssd1 vccd1 vccd1 _19624_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10473__C1 _10373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17457_ _16838_/X _19594_/Q _17457_/S vssd1 vssd1 vccd1 vccd1 _17458_/A sky130_fd_sc_hd__mux2_1
X_14669_ _14677_/A _15956_/B vssd1 vssd1 vccd1 vccd1 _14670_/A sky130_fd_sc_hd__and2_1
X_16408_ _16408_/A vssd1 vssd1 vccd1 vccd1 _19168_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15060__A _18456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17388_ _17388_/A vssd1 vssd1 vccd1 vccd1 _19563_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_164_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19506_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13962__A0 _18431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16339_ _16339_/A vssd1 vssd1 vccd1 vccd1 _19138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19127_ _19609_/CLK _19127_/D vssd1 vssd1 vccd1 vccd1 _19127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19058_ _19710_/CLK _19058_/D vssd1 vssd1 vccd1 vccd1 _19058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18009_ _18027_/A _18009_/B vssd1 vssd1 vccd1 vccd1 _18009_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_179_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19569_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13190__A1 _19664_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10623__S0 _10605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17208__A1 _12656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_102_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _18386_/CLK sky130_fd_sc_hd__clkbuf_16
X_09713_ _19527_/Q _19141_/Q _19591_/Q _18747_/Q _10257_/S _09542_/A vssd1 vssd1 vccd1
+ vccd1 _09714_/B sky130_fd_sc_hd__mux4_1
XFILLER_19_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17759__A2 _13399_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14690__A1 _14584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10926__S1 _10906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15235__A _16737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14690__B2 input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09644_ _09171_/A _09643_/X _10379_/A vssd1 vssd1 vccd1 vccd1 _09644_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09233__A _09854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09575_ _09732_/A vssd1 vssd1 vccd1 vccd1 _10182_/A sky130_fd_sc_hd__buf_2
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_117_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _18567_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_64_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13402__C1 _13401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10216__C1 _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13202__B _18625_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10350_ _18863_/Q _19321_/Q _10350_/S vssd1 vssd1 vccd1 vccd1 _10350_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10862__S0 _10614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09909__C1 _09231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10281_ _09735_/A _10278_/Y _10280_/Y _11119_/A vssd1 vssd1 vccd1 vccd1 _10281_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16005__S _16005_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12020_ _18363_/Q _18362_/Q _12020_/C vssd1 vssd1 vccd1 vccd1 _12075_/C sky130_fd_sc_hd__and3_1
XANTENNA__09924__A2 _09624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15844__S _15852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13971_ _14150_/A vssd1 vssd1 vccd1 vccd1 _13971_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14681__A1 _14578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11673__A _18343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15710_ _15721_/A vssd1 vssd1 vccd1 vccd1 _15719_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__14681__B2 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12922_ _17993_/A vssd1 vssd1 vccd1 vccd1 _12922_/X sky130_fd_sc_hd__buf_4
XFILLER_46_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16690_ _16722_/A vssd1 vssd1 vccd1 vccd1 _16703_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_47_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15641_ _18838_/Q _15558_/X _15647_/S vssd1 vssd1 vccd1 vccd1 _15642_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11392__B _11723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09143__A _09695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12853_ _18170_/A vssd1 vssd1 vccd1 vccd1 _12897_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16675__S _16687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _18395_/CLK _18360_/D vssd1 vssd1 vccd1 vccd1 _18360_/Q sky130_fd_sc_hd__dfxtp_2
X_11804_ _11804_/A vssd1 vssd1 vccd1 vccd1 _11804_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12444__A0 _11205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15572_ _18810_/Q _15570_/X _15584_/S vssd1 vssd1 vccd1 vccd1 _15573_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _18525_/Q _18524_/Q _18523_/Q _18522_/Q vssd1 vssd1 vccd1 vccd1 _12790_/C
+ sky130_fd_sc_hd__or4bb_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _19529_/Q _16731_/X _17313_/S vssd1 vssd1 vccd1 vccd1 _17312_/A sky130_fd_sc_hd__mux2_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14523_ _14577_/A vssd1 vssd1 vccd1 vccd1 _14551_/B sky130_fd_sc_hd__clkbuf_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18291_ _18298_/CLK _18291_/D vssd1 vssd1 vccd1 vccd1 _18291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _18578_/Q _14559_/A _11735_/S vssd1 vssd1 vccd1 vccd1 _11736_/C sky130_fd_sc_hd__mux2_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19798_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11612__S _15095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17242_ _19499_/Q _17241_/X _17245_/S vssd1 vssd1 vccd1 vccd1 _17243_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14454_ _18499_/Q _19737_/Q _14454_/S vssd1 vssd1 vccd1 vccd1 _14455_/A sky130_fd_sc_hd__mux2_1
X_11666_ _11749_/A vssd1 vssd1 vccd1 vccd1 _12411_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__14736__A2 _13163_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13405_ _19498_/Q _13203_/A _13115_/A _18379_/Q _13404_/X vssd1 vssd1 vccd1 vccd1
+ _13407_/A sky130_fd_sc_hd__a221o_1
XANTENNA__10207__C1 _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17173_ _17173_/A vssd1 vssd1 vccd1 vccd1 _19478_/D sky130_fd_sc_hd__clkbuf_1
X_10617_ _18761_/Q _18990_/Q _18921_/Q _19219_/Q _10614_/X _10616_/X vssd1 vssd1 vccd1
+ vccd1 _10618_/B sky130_fd_sc_hd__mux4_1
XFILLER_167_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14385_ _14883_/A _18505_/Q _14395_/S vssd1 vssd1 vccd1 vccd1 _14386_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14923__S _14923_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11597_ _12511_/A vssd1 vssd1 vccd1 vccd1 _11624_/A sky130_fd_sc_hd__clkinv_2
X_16124_ _16124_/A vssd1 vssd1 vccd1 vccd1 _19041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13336_ _13267_/X _13334_/X _13335_/X _13317_/X vssd1 vssd1 vccd1 vccd1 _18371_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_96_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19472_/CLK sky130_fd_sc_hd__clkbuf_16
X_10548_ _10548_/A vssd1 vssd1 vccd1 vccd1 _10548_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16055_ _16765_/A vssd1 vssd1 vccd1 vccd1 _16055_/X sky130_fd_sc_hd__clkbuf_1
X_13267_ _13354_/A vssd1 vssd1 vccd1 vccd1 _13267_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10479_ _19608_/Q _19446_/Q _18892_/Q _18662_/Q _09449_/A _09634_/A vssd1 vssd1 vccd1
+ vccd1 _10480_/B sky130_fd_sc_hd__mux4_2
XFILLER_170_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15006_ _14875_/X _15005_/X _14842_/X vssd1 vssd1 vccd1 vccd1 _15006_/X sky130_fd_sc_hd__o21a_1
XFILLER_130_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09318__A _09318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12218_ _12218_/A _12267_/C vssd1 vssd1 vccd1 vccd1 _12218_/X sky130_fd_sc_hd__or2_1
XFILLER_142_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13198_ _13365_/A vssd1 vssd1 vccd1 vccd1 _13438_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_111_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19814_ _19818_/CLK _19814_/D vssd1 vssd1 vccd1 vccd1 _19814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12149_ _18368_/Q vssd1 vssd1 vccd1 vccd1 _13316_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10081__S1 _10080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17535__A _17535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19745_ _19753_/CLK _19745_/D vssd1 vssd1 vccd1 vccd1 _19745_/Q sky130_fd_sc_hd__dfxtp_4
X_16957_ _16957_/A vssd1 vssd1 vccd1 vccd1 _19386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15908_ _15908_/A vssd1 vssd1 vccd1 vccd1 _18956_/D sky130_fd_sc_hd__clkbuf_1
X_19676_ _19682_/CLK _19676_/D vssd1 vssd1 vccd1 vccd1 _19676_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_34_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19397_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16888_ _16888_/A vssd1 vssd1 vccd1 vccd1 _19356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18627_ _19692_/CLK _18627_/D vssd1 vssd1 vccd1 vccd1 _18627_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15839_ _14867_/X _18926_/Q _15841_/S vssd1 vssd1 vccd1 vccd1 _15840_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10199__A _10212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13227__A2 _12665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09360_ _10132_/A vssd1 vssd1 vccd1 vccd1 _09880_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09988__A _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18558_ _18564_/CLK _18558_/D vssd1 vssd1 vccd1 vccd1 _18558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17509_ _17520_/A vssd1 vssd1 vccd1 vccd1 _17518_/S sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_49_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19721_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09291_ _18576_/Q _18531_/Q vssd1 vssd1 vccd1 vccd1 _09291_/X sky130_fd_sc_hd__and2_1
XFILLER_162_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18489_ _19079_/CLK _18489_/D vssd1 vssd1 vccd1 vccd1 _18489_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_162_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14727__A2 _14703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15929__S _15935_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput120 _12487_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[18] sky130_fd_sc_hd__buf_2
Xoutput131 _12502_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[28] sky130_fd_sc_hd__buf_2
Xoutput142 _12475_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[9] sky130_fd_sc_hd__buf_2
XFILLER_82_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput153 _17890_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[18] sky130_fd_sc_hd__buf_2
XFILLER_121_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09228__A _09708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput164 _17907_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[28] sky130_fd_sc_hd__buf_2
XFILLER_82_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput175 _17872_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[9] sky130_fd_sc_hd__buf_2
XANTENNA__09462__S0 _10350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11493__A _11513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09627_ _09430_/A _09607_/X _09623_/X _09625_/X _09626_/Y vssd1 vssd1 vccd1 vccd1
+ _12503_/A sky130_fd_sc_hd__o32a_4
XFILLER_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16495__S _16497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09898__A _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09558_ _10348_/S vssd1 vssd1 vccd1 vccd1 _10417_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_71_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15412__B _15412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09489_ _10770_/S vssd1 vssd1 vccd1 vccd1 _10788_/S sky130_fd_sc_hd__buf_2
XFILLER_169_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10988__B1 _19694_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11520_ _14566_/A _11628_/A _11665_/C _11520_/D vssd1 vssd1 vccd1 vccd1 _13527_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_12_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12729__A1 _17774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15839__S _15841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11451_ _11716_/A _11463_/B _11463_/C vssd1 vssd1 vccd1 vccd1 _14718_/B sky130_fd_sc_hd__and3_2
XFILLER_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10402_ _18831_/Q _19385_/Q _19547_/Q _18799_/Q _11112_/S _10384_/X vssd1 vssd1 vccd1
+ vccd1 _10403_/B sky130_fd_sc_hd__mux4_1
X_14170_ _14130_/A _14167_/X _14169_/Y _13950_/X vssd1 vssd1 vccd1 vccd1 _14170_/X
+ sky130_fd_sc_hd__a31o_1
X_11382_ _11369_/Y _11379_/X _11381_/X _18417_/Q vssd1 vssd1 vccd1 vccd1 _13532_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13121_ _13297_/A vssd1 vssd1 vccd1 vccd1 _13121_/X sky130_fd_sc_hd__buf_2
XANTENNA__11072__A2_N _12465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10333_ _09732_/A _10332_/X _09616_/A vssd1 vssd1 vccd1 vccd1 _10333_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_139_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input54_A io_ibus_inst[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ _13055_/A _13055_/C _13011_/X vssd1 vssd1 vccd1 vccd1 _13052_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09138__A _10969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10264_ _09215_/A _10255_/X _10259_/X _10263_/X _09134_/A vssd1 vssd1 vccd1 vccd1
+ _10264_/X sky130_fd_sc_hd__a311o_1
XFILLER_97_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12003_ _11991_/Y _11998_/Y _17878_/A _12002_/X vssd1 vssd1 vccd1 vccd1 _12003_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_105_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17860_ _17862_/A _17860_/B vssd1 vssd1 vccd1 vccd1 _17861_/A sky130_fd_sc_hd__or2_1
X_10195_ _10196_/A _12487_/A vssd1 vssd1 vccd1 vccd1 _10197_/A sky130_fd_sc_hd__and2_1
X_16811_ _16809_/X _19327_/Q _16823_/S vssd1 vssd1 vccd1 vccd1 _16812_/A sky130_fd_sc_hd__mux2_1
X_17791_ _17791_/A vssd1 vssd1 vccd1 vccd1 _19698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12499__A _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19530_ _19626_/CLK _19530_/D vssd1 vssd1 vccd1 vccd1 _19530_/Q sky130_fd_sc_hd__dfxtp_1
X_16742_ _16742_/A vssd1 vssd1 vccd1 vccd1 _19306_/D sky130_fd_sc_hd__clkbuf_1
X_13954_ _13743_/X _13756_/X _13966_/S vssd1 vssd1 vccd1 vccd1 _13954_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10511__S _10511_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12905_ _18034_/A vssd1 vssd1 vccd1 vccd1 _17999_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09530__B1 _09529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19461_ _19722_/CLK _19461_/D vssd1 vssd1 vccd1 vccd1 _19461_/Q sky130_fd_sc_hd__dfxtp_1
X_16673_ _16673_/A vssd1 vssd1 vccd1 vccd1 _16673_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13885_ _13764_/X _13768_/X _13888_/S vssd1 vssd1 vccd1 vccd1 _13885_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18412_ _19788_/CLK _18412_/D vssd1 vssd1 vccd1 vccd1 _18412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12836_ _18261_/Q vssd1 vssd1 vccd1 vccd1 _12840_/B sky130_fd_sc_hd__buf_2
X_15624_ _15624_/A vssd1 vssd1 vccd1 vccd1 _18830_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ _19620_/CLK _19392_/D vssd1 vssd1 vccd1 vccd1 _19392_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09601__A _10384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18343_ _19759_/CLK _18343_/D vssd1 vssd1 vccd1 vccd1 _18343_/Q sky130_fd_sc_hd__dfxtp_2
X_15555_ _15571_/A vssd1 vssd1 vccd1 vccd1 _15568_/S sky130_fd_sc_hd__buf_4
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12767_ _13324_/A _18643_/Q vssd1 vssd1 vccd1 vccd1 _12767_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10979__B1 _12463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13123__A _13123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14506_ _17862_/A _14506_/B vssd1 vssd1 vccd1 vccd1 _14507_/A sky130_fd_sc_hd__or2_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18274_ _18386_/CLK _18274_/D vssd1 vssd1 vccd1 vccd1 _18274_/Q sky130_fd_sc_hd__dfxtp_1
X_11718_ _15263_/A _11678_/B _11717_/X vssd1 vssd1 vccd1 vccd1 _11719_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__16137__C _16919_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15486_ _15486_/A vssd1 vssd1 vccd1 vccd1 _18784_/D sky130_fd_sc_hd__clkbuf_1
X_12698_ _12780_/S _12714_/B _18205_/A vssd1 vssd1 vccd1 vccd1 _13090_/S sky130_fd_sc_hd__o21a_1
XFILLER_174_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17225_ _18451_/Q _13364_/X _17235_/S vssd1 vssd1 vccd1 vccd1 _17225_/X sky130_fd_sc_hd__mux2_1
X_14437_ _18491_/Q _19729_/Q _14443_/S vssd1 vssd1 vccd1 vccd1 _14438_/A sky130_fd_sc_hd__mux2_1
X_11649_ _11697_/S vssd1 vssd1 vccd1 vccd1 _11840_/A sky130_fd_sc_hd__buf_2
Xinput11 io_dbus_rdata[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_4
Xinput22 io_dbus_rdata[29] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_2
XFILLER_30_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput33 io_dbus_valid vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_4
XFILLER_174_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput44 io_ibus_inst[19] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_2
X_17156_ _17156_/A vssd1 vssd1 vccd1 vccd1 _19473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput55 io_ibus_inst[29] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__buf_2
XANTENNA__10826__S0 _09152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14368_ _14368_/A vssd1 vssd1 vccd1 vccd1 _18467_/D sky130_fd_sc_hd__clkbuf_1
Xinput66 io_ibus_valid vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__buf_2
XFILLER_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16107_ _16106_/X _19036_/Q _16113_/S vssd1 vssd1 vccd1 vccd1 _16108_/A sky130_fd_sc_hd__mux2_1
X_13319_ _18369_/Q _13319_/B vssd1 vssd1 vccd1 vccd1 _13319_/X sky130_fd_sc_hd__or2_1
XFILLER_155_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17087_ _17087_/A vssd1 vssd1 vccd1 vccd1 _19444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14299_ _13927_/X _14296_/Y _14298_/X _13982_/X vssd1 vssd1 vccd1 vccd1 _14299_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_115_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16038_ _16038_/A vssd1 vssd1 vccd1 vccd1 _19014_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14889__A _16793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_12_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17989_ _18033_/A _17989_/B _17990_/B vssd1 vssd1 vccd1 vccd1 _19781_/D sky130_fd_sc_hd__nor3_1
XFILLER_38_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19728_ _19738_/CLK _19728_/D vssd1 vssd1 vccd1 vccd1 _19728_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19659_ _19659_/CLK _19659_/D vssd1 vssd1 vccd1 vccd1 _19659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09412_ _09412_/A vssd1 vssd1 vccd1 vccd1 _09616_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15070__A1 _18489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09343_ _11188_/S vssd1 vssd1 vccd1 vccd1 _09344_/A sky130_fd_sc_hd__buf_6
XANTENNA__09511__A _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09274_ _09274_/A vssd1 vssd1 vccd1 vccd1 _09275_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_138_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11631__B2 _19729_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10293__S1 _11113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17175__A _17245_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13439__A2 _13437_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10951_ _19600_/Q _19438_/Q _18884_/Q _18654_/Q _10631_/A _10726_/X vssd1 vssd1 vccd1
+ vccd1 _10951_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13670_ _12446_/B _12510_/B _13724_/B vssd1 vssd1 vccd1 vccd1 _13670_/X sky130_fd_sc_hd__mux2_1
X_10882_ _19245_/Q _19016_/Q _18947_/Q _19341_/Q _10724_/X _10726_/X vssd1 vssd1 vccd1
+ vccd1 _10883_/B sky130_fd_sc_hd__mux4_2
XANTENNA__15061__A1 _14958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12621_ _18322_/Q vssd1 vssd1 vccd1 vccd1 _13033_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16953__S _16953_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15340_ _16847_/B _17391_/B vssd1 vssd1 vccd1 vccd1 _15397_/A sky130_fd_sc_hd__nor2_4
XFILLER_40_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12552_ _19872_/Q _12525_/X _12528_/X _19840_/Q _12551_/X vssd1 vssd1 vccd1 vccd1
+ _12552_/X sky130_fd_sc_hd__a221o_1
XFILLER_106_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11503_ _14580_/A _18578_/Q vssd1 vssd1 vccd1 vccd1 _11519_/D sky130_fd_sc_hd__or2_1
XFILLER_129_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15271_ _15271_/A vssd1 vssd1 vccd1 vccd1 _18689_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12483_ _12483_/A _12483_/B vssd1 vssd1 vccd1 vccd1 _12483_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17010_ _19410_/Q _16664_/X _17014_/S vssd1 vssd1 vccd1 vccd1 _17011_/A sky130_fd_sc_hd__mux2_1
X_14222_ _18447_/Q _11460_/A _14211_/Y _14221_/X vssd1 vssd1 vccd1 vccd1 _18447_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_172_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11434_ _18553_/Q _18552_/Q vssd1 vssd1 vccd1 vccd1 _11434_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14153_ _13978_/X _14155_/B _13797_/A _14152_/X vssd1 vssd1 vccd1 vccd1 _14153_/X
+ sky130_fd_sc_hd__o211a_1
X_11365_ _11365_/A _11365_/B _11528_/B vssd1 vssd1 vccd1 vccd1 _11365_/X sky130_fd_sc_hd__or3_1
XFILLER_164_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13104_ input70/X _13104_/B vssd1 vssd1 vccd1 vccd1 _13104_/X sky130_fd_sc_hd__or2_1
XFILLER_125_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10316_ _09172_/A _10315_/X _09184_/A vssd1 vssd1 vccd1 vccd1 _10316_/X sky130_fd_sc_hd__a21o_1
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14084_ _18437_/Q _11460_/X _14083_/X vssd1 vssd1 vccd1 vccd1 _18437_/D sky130_fd_sc_hd__o21a_1
X_18961_ _19452_/CLK _18961_/D vssd1 vssd1 vccd1 vccd1 _18961_/Q sky130_fd_sc_hd__dfxtp_1
X_11296_ _11585_/A _11501_/B _11296_/C _11468_/C vssd1 vssd1 vccd1 vccd1 _11564_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_106_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17912_ _19759_/Q _12186_/A _12454_/X _12456_/X _17895_/X vssd1 vssd1 vccd1 vccd1
+ _19759_/D sky130_fd_sc_hd__o221a_1
XFILLER_152_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13035_ _18322_/Q _18324_/Q _18323_/Q _13035_/D vssd1 vssd1 vccd1 vccd1 _13047_/D
+ sky130_fd_sc_hd__and4_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10247_ _19420_/Q _19196_/Q _19713_/Q _19164_/Q _11110_/S _09483_/X vssd1 vssd1 vccd1
+ vccd1 _10247_/X sky130_fd_sc_hd__mux4_1
X_18892_ _19608_/CLK _18892_/D vssd1 vssd1 vccd1 vccd1 _18892_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_186_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17843_ _15223_/X _19722_/Q _17849_/S vssd1 vssd1 vccd1 vccd1 _17844_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10178_ _19647_/Q _19064_/Q _19101_/Q _18707_/Q _09721_/X _09610_/X vssd1 vssd1 vccd1
+ vccd1 _10178_/X sky130_fd_sc_hd__mux4_1
XANTENNA__14627__A1 _18563_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17774_ _17774_/A _17774_/B vssd1 vssd1 vccd1 vccd1 _19691_/D sky130_fd_sc_hd__nor2_2
X_14986_ _16819_/A vssd1 vssd1 vccd1 vccd1 _14986_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19513_ _19513_/CLK _19513_/D vssd1 vssd1 vccd1 vccd1 _19513_/Q sky130_fd_sc_hd__dfxtp_1
X_16725_ _16725_/A vssd1 vssd1 vccd1 vccd1 _16725_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13937_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13937_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19444_ _19444_/CLK _19444_/D vssd1 vssd1 vccd1 vccd1 _19444_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11861__A1 _19735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16656_ _16656_/A vssd1 vssd1 vccd1 vccd1 _19279_/D sky130_fd_sc_hd__clkbuf_1
X_13868_ _13868_/A _13868_/B vssd1 vssd1 vccd1 vccd1 _13868_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15052__A1 _14744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12819_ _12821_/B _12821_/C _12818_/Y vssd1 vssd1 vccd1 vccd1 _18255_/D sky130_fd_sc_hd__o21a_1
X_15607_ _15607_/A vssd1 vssd1 vccd1 vccd1 _18822_/D sky130_fd_sc_hd__clkbuf_1
X_19375_ _19537_/CLK _19375_/D vssd1 vssd1 vccd1 vccd1 _19375_/Q sky130_fd_sc_hd__dfxtp_1
X_13799_ _14212_/A _13877_/S vssd1 vssd1 vccd1 vccd1 _13799_/Y sky130_fd_sc_hd__nand2_1
X_16587_ _19249_/Q vssd1 vssd1 vccd1 vccd1 _16588_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16863__S _16869_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18326_ _19822_/CLK _18326_/D vssd1 vssd1 vccd1 vccd1 _18326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15538_ _16793_/A vssd1 vssd1 vccd1 vccd1 _15538_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16001__A0 _14918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10196__B _12487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15479__S _15481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18257_ _19855_/CLK _18257_/D vssd1 vssd1 vccd1 vccd1 _18257_/Q sky130_fd_sc_hd__dfxtp_1
X_15469_ _15469_/A vssd1 vssd1 vccd1 vccd1 _18776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17208_ _18446_/Q _12656_/B _17218_/S vssd1 vssd1 vccd1 vccd1 _17208_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18188_ _19850_/Q _18191_/C _18170_/X vssd1 vssd1 vccd1 vccd1 _18188_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09665__S0 _10328_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17139_ _17226_/A vssd1 vssd1 vccd1 vccd1 _17245_/S sky130_fd_sc_hd__buf_2
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10275__S1 _10239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09961_ _19425_/Q _19201_/Q _19718_/Q _19169_/Q _09803_/A _09936_/X vssd1 vssd1 vccd1
+ vccd1 _09961_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09968__S1 _09936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09892_ _09892_/A vssd1 vssd1 vccd1 vccd1 _09892_/X sky130_fd_sc_hd__buf_2
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09506__A _10400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15942__S _15946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09326_ _10524_/A vssd1 vssd1 vccd1 vccd1 _10496_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15389__S _15395_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13698__A _13702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09257_ _18530_/Q vssd1 vssd1 vccd1 vccd1 _16138_/A sky130_fd_sc_hd__clkinv_2
XFILLER_166_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16074__A _16784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13357__A1 _19684_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09188_ _09788_/A vssd1 vssd1 vccd1 vccd1 _09237_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14306__A0 _18454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ _11150_/A vssd1 vssd1 vccd1 vccd1 _11151_/C sky130_fd_sc_hd__inv_2
X_10101_ _10098_/X _12489_/C vssd1 vssd1 vccd1 vccd1 _10102_/B sky130_fd_sc_hd__and2b_1
XFILLER_136_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11081_ _11081_/A vssd1 vssd1 vccd1 vccd1 _11081_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09959__S1 _09869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14322__A _14324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ _09936_/X _10032_/B vssd1 vssd1 vccd1 vccd1 _10032_/X sky130_fd_sc_hd__and2b_1
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15852__S _15852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11157__S _11157_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14840_ _18469_/Q _14840_/B vssd1 vssd1 vccd1 vccd1 _14861_/C sky130_fd_sc_hd__and2_1
XFILLER_64_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14771_ _16657_/A vssd1 vssd1 vccd1 vccd1 _16761_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input17_A io_dbus_rdata[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ _11901_/C _12093_/D _17878_/A vssd1 vssd1 vccd1 vccd1 _11985_/A sky130_fd_sc_hd__a21oi_1
XFILLER_57_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16510_ _19213_/Q _15497_/X _16514_/S vssd1 vssd1 vccd1 vccd1 _16511_/A sky130_fd_sc_hd__mux2_1
X_13722_ _13747_/S _13714_/X _13719_/X _11624_/A _13721_/X vssd1 vssd1 vccd1 vccd1
+ _13722_/X sky130_fd_sc_hd__a221o_1
X_10934_ _18589_/Q _19278_/Q _10934_/S vssd1 vssd1 vccd1 vccd1 _10934_/X sky130_fd_sc_hd__mux2_1
X_17490_ _19608_/Q _16677_/X _17496_/S vssd1 vssd1 vccd1 vccd1 _17491_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09151__A _11028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13653_ _13653_/A vssd1 vssd1 vccd1 vccd1 _14034_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_16441_ _16441_/A vssd1 vssd1 vccd1 vccd1 _19182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ _18758_/Q _18987_/Q _18918_/Q _19216_/Q _09152_/A _10740_/A vssd1 vssd1 vccd1
+ vccd1 _10866_/B sky130_fd_sc_hd__mux4_1
XFILLER_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12604_ _12604_/A vssd1 vssd1 vccd1 vccd1 _12604_/X sky130_fd_sc_hd__clkbuf_2
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14793__A0 _14792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19160_ _19707_/CLK _19160_/D vssd1 vssd1 vccd1 vccd1 _19160_/Q sky130_fd_sc_hd__dfxtp_1
X_16372_ _19152_/Q _15506_/X _16380_/S vssd1 vssd1 vccd1 vccd1 _16373_/A sky130_fd_sc_hd__mux2_1
X_13584_ _13584_/A _13584_/B _13584_/C _13584_/D vssd1 vssd1 vccd1 vccd1 _13585_/D
+ sky130_fd_sc_hd__or4_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ _19407_/Q _19183_/Q _19700_/Q _19151_/Q _10934_/S _10713_/A vssd1 vssd1 vccd1
+ vccd1 _10797_/B sky130_fd_sc_hd__mux4_1
XANTENNA__18183__B _19847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15323_ _15323_/A vssd1 vssd1 vccd1 vccd1 _18713_/D sky130_fd_sc_hd__clkbuf_1
X_18111_ _18120_/A _18111_/B _18111_/C vssd1 vssd1 vccd1 vccd1 _19824_/D sky130_fd_sc_hd__nor3_1
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ _12751_/C _12566_/A _12670_/C vssd1 vssd1 vccd1 vccd1 _12587_/A sky130_fd_sc_hd__and3b_1
XFILLER_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19091_ _19638_/CLK _19091_/D vssd1 vssd1 vccd1 vccd1 _19091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18042_ _18085_/A vssd1 vssd1 vccd1 vccd1 _18077_/A sky130_fd_sc_hd__buf_2
X_15254_ _17762_/S _15254_/B vssd1 vssd1 vccd1 vccd1 _15255_/B sky130_fd_sc_hd__nor2_2
XFILLER_9_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12466_ _12466_/A _12466_/B vssd1 vssd1 vccd1 vccd1 _12467_/A sky130_fd_sc_hd__and2_1
XFILLER_144_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14216__B _14216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14205_ _13788_/A _14202_/X _14204_/Y _13894_/A vssd1 vssd1 vccd1 vccd1 _14205_/X
+ sky130_fd_sc_hd__a31o_1
X_11417_ _12533_/A _12533_/B _11821_/A _12540_/A vssd1 vssd1 vccd1 vccd1 _11419_/C
+ sky130_fd_sc_hd__or4b_2
X_15185_ _18665_/Q _15184_/X _15185_/S vssd1 vssd1 vccd1 vccd1 _15186_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12017__A _19672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12397_ _12419_/A _12397_/B vssd1 vssd1 vccd1 vccd1 _14310_/B sky130_fd_sc_hd__nand2_2
XANTENNA__16712__A _16712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14136_ _13753_/X _13994_/Y _14135_/Y _14086_/S vssd1 vssd1 vccd1 vccd1 _14136_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_output85_A _12185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11348_ _11372_/A _11343_/X _11345_/Y _11347_/Y vssd1 vssd1 vccd1 vccd1 _11587_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10582__A1 _10238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10881__A1_N _12465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17019__S _17025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18944_ _19804_/CLK _18944_/D vssd1 vssd1 vccd1 vccd1 _18944_/Q sky130_fd_sc_hd__dfxtp_1
X_14067_ _14054_/X _14056_/X _14066_/X _13784_/X vssd1 vssd1 vccd1 vccd1 _14067_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11279_ _11284_/C _11219_/X _11278_/Y vssd1 vssd1 vccd1 vccd1 _11279_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_140_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13018_ _13026_/D vssd1 vssd1 vccd1 vccd1 _13024_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18875_ _19397_/CLK _18875_/D vssd1 vssd1 vccd1 vccd1 _18875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17826_ _17826_/A vssd1 vssd1 vccd1 vccd1 _19714_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14076__A2 _14074_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17757_ _18486_/Q _17757_/B vssd1 vssd1 vccd1 vccd1 _17757_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14969_ _14969_/A _14969_/B _14978_/B vssd1 vssd1 vccd1 vccd1 _14969_/X sky130_fd_sc_hd__or3_1
XFILLER_75_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16708_ _16708_/A vssd1 vssd1 vccd1 vccd1 _19295_/D sky130_fd_sc_hd__clkbuf_1
X_17688_ _19674_/Q _17686_/X _17718_/S vssd1 vssd1 vccd1 vccd1 _17689_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11834__B2 _10810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15025__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19427_ _19427_/CLK _19427_/D vssd1 vssd1 vccd1 vccd1 _19427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16639_ _16639_/A vssd1 vssd1 vccd1 vccd1 _16639_/X sky130_fd_sc_hd__buf_2
XFILLER_149_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09996__A _09996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19358_ _19648_/CLK _19358_/D vssd1 vssd1 vccd1 vccd1 _19358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09111_ _18567_/Q vssd1 vssd1 vccd1 vccd1 _11365_/B sky130_fd_sc_hd__inv_2
X_18309_ _18329_/CLK _18309_/D vssd1 vssd1 vccd1 vccd1 _18309_/Q sky130_fd_sc_hd__dfxtp_1
X_19289_ _19513_/CLK _19289_/D vssd1 vssd1 vccd1 vccd1 _19289_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13339__A1 _19681_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13545__A_N _13578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14126__B _14126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14839__A1 _12711_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09944_ _09944_/A _09944_/B vssd1 vssd1 vccd1 vccd1 _09944_/X sky130_fd_sc_hd__or2_1
XANTENNA__10670__A _10813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09875_ _09875_/A _09875_/B vssd1 vssd1 vccd1 vccd1 _09875_/Y sky130_fd_sc_hd__nand2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input9_A io_dbus_rdata[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12078__B2 _12485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17599__S _17601_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_134_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10650_ _18594_/Q _19283_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _10651_/B sky130_fd_sc_hd__mux2_1
XFILLER_70_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09877__S0 _09803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09309_ _09309_/A vssd1 vssd1 vccd1 vccd1 _09309_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10581_ _18595_/Q _19284_/Q _10581_/S vssd1 vssd1 vccd1 vccd1 _10581_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16008__S _16016_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12320_ _18375_/Q _13352_/A _12320_/C vssd1 vssd1 vccd1 vccd1 _12341_/B sky130_fd_sc_hd__and3_1
XFILLER_108_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12251_ _18372_/Q _12272_/C vssd1 vssd1 vccd1 vccd1 _12251_/X sky130_fd_sc_hd__and2_1
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11202_ _11202_/A _12504_/A vssd1 vssd1 vccd1 vccd1 _11203_/B sky130_fd_sc_hd__nor2_1
XFILLER_134_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12182_ _12182_/A _12182_/B vssd1 vssd1 vccd1 vccd1 _12185_/A sky130_fd_sc_hd__nor2_2
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11761__B1 _11716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11133_ _11130_/Y _10462_/A _11131_/A vssd1 vssd1 vccd1 vccd1 _11133_/Y sky130_fd_sc_hd__a21oi_1
X_16990_ _16844_/X _19402_/Q _16990_/S vssd1 vssd1 vccd1 vccd1 _16991_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13502__A1 _13376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15941_ _15941_/A vssd1 vssd1 vccd1 vccd1 _18971_/D sky130_fd_sc_hd__clkbuf_1
X_11064_ _18817_/Q _19371_/Q _19533_/Q _18785_/Q _10805_/A _10725_/A vssd1 vssd1 vccd1
+ vccd1 _11065_/B sky130_fd_sc_hd__mux4_1
XFILLER_1_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10316__A1 _09172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_59_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16678__S _16687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12710__C1 _12709_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10015_ _18774_/Q _19003_/Q _18934_/Q _19232_/Q _10076_/S _09979_/A vssd1 vssd1 vccd1
+ vccd1 _10016_/B sky130_fd_sc_hd__mux4_1
XFILLER_88_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17244__A2 _17628_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18660_ _19444_/CLK _18660_/D vssd1 vssd1 vccd1 vccd1 _18660_/Q sky130_fd_sc_hd__dfxtp_1
X_15872_ _15044_/X _18941_/Q _15874_/S vssd1 vssd1 vccd1 vccd1 _15873_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14058__A2 _14057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17611_ _19082_/Q _17611_/B vssd1 vssd1 vccd1 vccd1 _17611_/Y sky130_fd_sc_hd__nand2_1
X_14823_ _14823_/A vssd1 vssd1 vccd1 vccd1 _18595_/D sky130_fd_sc_hd__clkbuf_1
X_18591_ _19506_/CLK _18591_/D vssd1 vssd1 vccd1 vccd1 _18591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17542_ _19631_/Q _16752_/A _17546_/S vssd1 vssd1 vccd1 vccd1 _17543_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14754_ _14753_/X _18589_/Q _14762_/S vssd1 vssd1 vccd1 vccd1 _14755_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11966_ _12024_/A _11966_/B vssd1 vssd1 vccd1 vccd1 _12026_/A sky130_fd_sc_hd__or2_1
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ _13702_/A _11733_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13706_/B sky130_fd_sc_hd__o21ai_2
X_10917_ _19695_/Q _10917_/B _10917_/C vssd1 vssd1 vccd1 vccd1 _10917_/X sky130_fd_sc_hd__or3_1
X_14685_ _14694_/A _14685_/B vssd1 vssd1 vccd1 vccd1 _14686_/A sky130_fd_sc_hd__and2_1
X_17473_ _17473_/A vssd1 vssd1 vccd1 vccd1 _19600_/D sky130_fd_sc_hd__clkbuf_1
X_11897_ _11922_/A _13614_/A vssd1 vssd1 vccd1 vccd1 _11899_/A sky130_fd_sc_hd__xor2_4
XFILLER_60_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17302__S _17302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19212_ _19696_/CLK _19212_/D vssd1 vssd1 vccd1 vccd1 _19212_/Q sky130_fd_sc_hd__dfxtp_1
X_13636_ _13658_/A _12282_/A _13685_/S vssd1 vssd1 vccd1 vccd1 _13636_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16424_ _19176_/Q _15583_/X _16424_/S vssd1 vssd1 vccd1 vccd1 _16425_/A sky130_fd_sc_hd__mux2_1
X_10848_ _10899_/A _10848_/B vssd1 vssd1 vccd1 vccd1 _10848_/X sky130_fd_sc_hd__or2_1
XFILLER_44_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19143_ _19657_/CLK _19143_/D vssd1 vssd1 vccd1 vccd1 _19143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17704__A0 _12617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13567_ _13567_/A vssd1 vssd1 vccd1 vccd1 _13720_/A sky130_fd_sc_hd__clkbuf_4
X_16355_ _16134_/X _19146_/Q _16355_/S vssd1 vssd1 vccd1 vccd1 _16356_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10478__S1 _09635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10779_ _10803_/A _10776_/X _10778_/X _10728_/X vssd1 vssd1 vccd1 vccd1 _10780_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14227__A _14227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12518_ _12518_/A vssd1 vssd1 vccd1 vccd1 _12518_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15306_ _15306_/A vssd1 vssd1 vccd1 vccd1 _18705_/D sky130_fd_sc_hd__clkbuf_1
X_19074_ _19657_/CLK _19074_/D vssd1 vssd1 vccd1 vccd1 _19074_/Q sky130_fd_sc_hd__dfxtp_1
X_16286_ _16342_/A vssd1 vssd1 vccd1 vccd1 _16355_/S sky130_fd_sc_hd__buf_6
X_13498_ _13498_/A vssd1 vssd1 vccd1 vccd1 _18407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18025_ _18033_/A _18025_/B _18025_/C vssd1 vssd1 vccd1 vccd1 _19794_/D sky130_fd_sc_hd__nor3_1
XFILLER_60_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15237_ _15237_/A vssd1 vssd1 vccd1 vccd1 _18681_/D sky130_fd_sc_hd__clkbuf_1
X_12449_ _13590_/S _12449_/B vssd1 vssd1 vccd1 vccd1 _12450_/B sky130_fd_sc_hd__xnor2_2
XFILLER_160_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15168_ _16670_/A vssd1 vssd1 vccd1 vccd1 _15168_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_154_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14119_ _14119_/A vssd1 vssd1 vccd1 vccd1 _18439_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15058__A _18488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15099_ _18625_/Q _13566_/X _15097_/X _11075_/A vssd1 vssd1 vccd1 vccd1 _18625_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18927_ _19223_/CLK _18927_/D vssd1 vssd1 vccd1 vccd1 _18927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09660_ _18844_/Q _19398_/Q _19560_/Q _18812_/Q _09600_/A _09603_/A vssd1 vssd1 vccd1
+ vccd1 _09661_/B sky130_fd_sc_hd__mux4_1
X_18858_ _19541_/CLK _18858_/D vssd1 vssd1 vccd1 vccd1 _18858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15246__A1 _11820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17809_ _17809_/A vssd1 vssd1 vccd1 vccd1 _19706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09591_ _10242_/S vssd1 vssd1 vccd1 vccd1 _09675_/S sky130_fd_sc_hd__buf_4
X_18789_ _19537_/CLK _18789_/D vssd1 vssd1 vccd1 vccd1 _18789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10166__S0 _10200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14757__A0 _10810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09859__S0 _09163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12232__A1 _10003_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10469__S1 _09635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17171__A1 _13245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13976__A _13984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10641__S1 _10634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09927_ _09927_/A vssd1 vssd1 vccd1 vccd1 _09927_/X sky130_fd_sc_hd__buf_4
XFILLER_59_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_60_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09858_ _09905_/A _09858_/B vssd1 vssd1 vccd1 vccd1 _09858_/X sky130_fd_sc_hd__or2_1
XANTENNA__14600__A _14612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _19525_/Q _19139_/Q _19589_/Q _18745_/Q _09760_/X _09841_/A vssd1 vssd1 vccd1
+ vccd1 _09790_/B sky130_fd_sc_hd__mux4_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _18356_/Q _11820_/B vssd1 vssd1 vccd1 vccd1 _11826_/A sky130_fd_sc_hd__xnor2_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _12119_/S _11751_/B vssd1 vssd1 vccd1 vccd1 _11751_/X sky130_fd_sc_hd__or2_1
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16527__A _16573_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17122__S _17130_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10702_ _18824_/Q _19378_/Q _19540_/Q _18792_/Q _10770_/S _09512_/A vssd1 vssd1 vccd1
+ vccd1 _10702_/X sky130_fd_sc_hd__mux4_2
XFILLER_53_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _18506_/Q _12095_/A _14476_/S vssd1 vssd1 vccd1 vccd1 _14471_/A sky130_fd_sc_hd__mux2_1
X_11682_ _11678_/X _11679_/Y _17241_/S vssd1 vssd1 vccd1 vccd1 _11682_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_41_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _19822_/Q _12665_/X _12602_/X _18333_/Q _13420_/X vssd1 vssd1 vccd1 vccd1
+ _13422_/B sky130_fd_sc_hd__a221o_4
XANTENNA__12223__A1 _17730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10633_ _10785_/A vssd1 vssd1 vccd1 vccd1 _10634_/A sky130_fd_sc_hd__buf_2
XFILLER_167_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12493__C _12493_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16140_ _16196_/A vssd1 vssd1 vccd1 vccd1 _16209_/S sky130_fd_sc_hd__buf_6
XANTENNA__12774__A2 _13130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13352_ _13352_/A _13352_/B vssd1 vssd1 vccd1 vccd1 _13352_/X sky130_fd_sc_hd__or2_1
XFILLER_10_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10564_ _19412_/Q _19188_/Q _19705_/Q _19156_/Q _10466_/S _09141_/A vssd1 vssd1 vccd1
+ vccd1 _10564_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12303_ _12323_/A _12303_/B vssd1 vssd1 vccd1 vccd1 _14265_/A sky130_fd_sc_hd__nand2_4
XFILLER_154_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16071_ _16781_/A vssd1 vssd1 vccd1 vccd1 _16071_/X sky130_fd_sc_hd__clkbuf_2
X_13283_ _13267_/X _13279_/X _13280_/X _13282_/X vssd1 vssd1 vccd1 vccd1 _18363_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10495_ _19512_/Q _19126_/Q _19576_/Q _18732_/Q _10242_/S _10239_/A vssd1 vssd1 vccd1
+ vccd1 _10496_/B sky130_fd_sc_hd__mux4_2
XFILLER_5_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15022_ _16829_/A vssd1 vssd1 vccd1 vccd1 _15022_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12234_ _12234_/A vssd1 vssd1 vccd1 vccd1 _12240_/A sky130_fd_sc_hd__inv_2
XFILLER_5_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19830_ _19833_/CLK _19830_/D vssd1 vssd1 vccd1 vccd1 _19830_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_122_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17792__S _17794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12165_ _12163_/Y _12164_/X _12165_/S vssd1 vssd1 vccd1 vccd1 _12165_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11116_ _10447_/A _11111_/X _11113_/Y _11115_/Y vssd1 vssd1 vccd1 vccd1 _11116_/X
+ sky130_fd_sc_hd__a31o_1
X_19761_ _19822_/CLK _19761_/D vssd1 vssd1 vccd1 vccd1 _19761_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_123_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16973_ _16819_/X _19394_/Q _16975_/S vssd1 vssd1 vccd1 vccd1 _16974_/A sky130_fd_sc_hd__mux2_1
X_12096_ _12408_/A _12096_/B vssd1 vssd1 vccd1 vccd1 _12096_/X sky130_fd_sc_hd__and2b_1
XFILLER_111_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18712_ _19718_/CLK _18712_/D vssd1 vssd1 vccd1 vccd1 _18712_/Q sky130_fd_sc_hd__dfxtp_1
X_15924_ _14940_/X _18964_/Q _15924_/S vssd1 vssd1 vccd1 vccd1 _15925_/A sky130_fd_sc_hd__mux2_1
X_11047_ _10857_/X _11035_/X _11044_/X _11046_/Y vssd1 vssd1 vccd1 vccd1 _11047_/X
+ sky130_fd_sc_hd__o31a_1
X_19692_ _19692_/CLK _19692_/D vssd1 vssd1 vccd1 vccd1 _19692_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16201__S _16205_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10396__S0 _09673_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 io_dbus_rdata[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_2
XFILLER_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18643_ _19628_/CLK _18643_/D vssd1 vssd1 vccd1 vccd1 _18643_/Q sky130_fd_sc_hd__dfxtp_1
X_15855_ _14951_/X _18933_/Q _15863_/S vssd1 vssd1 vccd1 vccd1 _15856_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10170__C1 _09249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14806_ _11542_/X _14800_/X _14805_/X vssd1 vssd1 vccd1 vccd1 _16667_/A sky130_fd_sc_hd__o21a_2
XFILLER_149_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18574_ _18618_/CLK _18574_/D vssd1 vssd1 vccd1 vccd1 _18574_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15786_ _15786_/A vssd1 vssd1 vccd1 vccd1 _18902_/D sky130_fd_sc_hd__clkbuf_1
X_12998_ _18312_/Q _12994_/C _12997_/Y vssd1 vssd1 vccd1 vccd1 _18312_/D sky130_fd_sc_hd__o21a_1
XFILLER_92_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17525_ _19624_/Q _16728_/X _17529_/S vssd1 vssd1 vccd1 vccd1 _17526_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14737_ _14737_/A _14743_/A vssd1 vssd1 vccd1 vccd1 _14737_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__09863__C1 _09249_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12965__A _18225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ _18501_/Q _12259_/B _12259_/C vssd1 vssd1 vccd1 vccd1 _11949_/X sky130_fd_sc_hd__or3_2
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17032__S _17036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15341__A _15397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17456_ _17456_/A vssd1 vssd1 vccd1 vccd1 _19593_/D sky130_fd_sc_hd__clkbuf_1
X_14668_ _14568_/A _12660_/A _14640_/A input48/X vssd1 vssd1 vccd1 vccd1 _15956_/B
+ sky130_fd_sc_hd__a22o_1
X_16407_ _19168_/Q _15558_/X _16413_/S vssd1 vssd1 vccd1 vccd1 _16408_/A sky130_fd_sc_hd__mux2_1
X_13619_ _13616_/X _13618_/X _13758_/S vssd1 vssd1 vccd1 vccd1 _13619_/X sky130_fd_sc_hd__mux2_1
X_17387_ _16841_/X _19563_/Q _17389_/S vssd1 vssd1 vccd1 vccd1 _17388_/A sky130_fd_sc_hd__mux2_1
X_14599_ _11297_/B _14597_/X _14593_/X _14598_/Y vssd1 vssd1 vccd1 vccd1 _14600_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_158_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19126_ _19608_/CLK _19126_/D vssd1 vssd1 vccd1 vccd1 _19126_/Q sky130_fd_sc_hd__dfxtp_1
X_16338_ _16109_/X _19138_/Q _16340_/S vssd1 vssd1 vccd1 vccd1 _16339_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19057_ _19640_/CLK _19057_/D vssd1 vssd1 vccd1 vccd1 _19057_/Q sky130_fd_sc_hd__dfxtp_1
X_16269_ _16269_/A vssd1 vssd1 vccd1 vccd1 _19107_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16900__A1 _16715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18008_ _19788_/Q _18011_/C vssd1 vssd1 vccd1 vccd1 _18009_/B sky130_fd_sc_hd__and2_1
XANTENNA__14911__A0 _18443_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10528__B2 _18436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10623__S1 _10366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12205__A _14216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09712_ _09712_/A _09712_/B vssd1 vssd1 vccd1 vccd1 _09712_/X sky130_fd_sc_hd__or2_1
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09514__A _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09643_ _18876_/Q _19334_/Q _09643_/S vssd1 vssd1 vccd1 vccd1 _09643_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10161__C1 _09135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15950__S _15950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09574_ _09276_/A _09564_/X _09573_/X _09283_/A _18455_/Q vssd1 vssd1 vccd1 vccd1
+ _11200_/A sky130_fd_sc_hd__a32o_4
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12594__B _12594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10395__A _10395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10862__S1 _10616_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13705__A1 _13702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10280_ _10280_/A _10280_/B vssd1 vssd1 vccd1 vccd1 _10280_/Y sky130_fd_sc_hd__nand2_1
XFILLER_152_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12115__A _14163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_0_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19609_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17117__S _17119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16021__S _16027_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13970_ _13967_/X _13969_/X _13970_/S vssd1 vssd1 vccd1 vccd1 _13970_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10378__S0 _09448_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12921_ _18034_/A vssd1 vssd1 vccd1 vccd1 _17993_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16956__S _16964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17080__A0 _16765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15640_ _15640_/A vssd1 vssd1 vccd1 vccd1 _18837_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _18034_/A vssd1 vssd1 vccd1 vccd1 _18170_/A sky130_fd_sc_hd__buf_4
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _11803_/A _11803_/B vssd1 vssd1 vccd1 vccd1 _11804_/A sky130_fd_sc_hd__and2_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15571_ _15571_/A vssd1 vssd1 vccd1 vccd1 _15584_/S sky130_fd_sc_hd__clkbuf_8
X_12783_ _18533_/Q _14716_/A _15134_/A vssd1 vssd1 vccd1 vccd1 _16847_/A sky130_fd_sc_hd__or3_4
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10455__B1 _09314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _17310_/A vssd1 vssd1 vccd1 vccd1 _19528_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ _14572_/B vssd1 vssd1 vccd1 vccd1 _14522_/X sky130_fd_sc_hd__clkbuf_2
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ _18573_/Q vssd1 vssd1 vccd1 vccd1 _14559_/A sky130_fd_sc_hd__clkbuf_4
X_18290_ _18298_/CLK _18290_/D vssd1 vssd1 vccd1 vccd1 _18290_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _18456_/Q _13423_/X _17241_/S vssd1 vssd1 vccd1 vccd1 _17241_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14197__A1 _12163_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14453_ _14453_/A vssd1 vssd1 vccd1 vccd1 _18498_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16691__S _16703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11665_ _19730_/Q _11665_/B _11665_/C _11665_/D vssd1 vssd1 vccd1 vccd1 _11665_/X
+ sky130_fd_sc_hd__or4_2
X_13404_ _18296_/Q _13404_/B vssd1 vssd1 vccd1 vccd1 _13404_/X sky130_fd_sc_hd__and2_1
X_10616_ _10906_/A vssd1 vssd1 vccd1 vccd1 _10616_/X sky130_fd_sc_hd__buf_4
XFILLER_168_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17172_ _19478_/Q _17171_/X _17172_/S vssd1 vssd1 vccd1 vccd1 _17173_/A sky130_fd_sc_hd__mux2_1
X_14384_ _14384_/A vssd1 vssd1 vccd1 vccd1 _14395_/S sky130_fd_sc_hd__clkbuf_2
X_11596_ _13625_/A _12510_/B vssd1 vssd1 vccd1 vccd1 _12511_/A sky130_fd_sc_hd__and2_2
XANTENNA__18191__B _19850_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10758__B2 _18432_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13335_ _18371_/Q _13352_/B vssd1 vssd1 vccd1 vccd1 _13335_/X sky130_fd_sc_hd__or2_1
XFILLER_127_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16123_ _16122_/X _19041_/Q _16129_/S vssd1 vssd1 vccd1 vccd1 _16124_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17088__A _17134_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10547_ _10813_/A vssd1 vssd1 vccd1 vccd1 _10548_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_157_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13266_ _12727_/X _13118_/X _13265_/X _13232_/X vssd1 vssd1 vccd1 vccd1 _18362_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16054_ _16054_/A vssd1 vssd1 vccd1 vccd1 _19019_/D sky130_fd_sc_hd__clkbuf_1
X_10478_ _18828_/Q _19382_/Q _19544_/Q _18796_/Q _09447_/A _09635_/A vssd1 vssd1 vccd1
+ vccd1 _10478_/X sky130_fd_sc_hd__mux4_1
XFILLER_142_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14224__B _14227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12217_ _19749_/Q _12217_/B vssd1 vssd1 vccd1 vccd1 _12267_/C sky130_fd_sc_hd__and2_1
X_15005_ _18451_/Q _13363_/B _15071_/S vssd1 vssd1 vccd1 vccd1 _15005_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13197_ _13121_/X _13187_/Y _13196_/X _13135_/X _18624_/Q vssd1 vssd1 vccd1 vccd1
+ _13197_/X sky130_fd_sc_hd__a32o_4
XFILLER_29_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11183__A1 _09616_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__A0 _11199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19813_ _19818_/CLK _19813_/D vssd1 vssd1 vccd1 vccd1 _19813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12148_ _12098_/B _12146_/X _12147_/Y vssd1 vssd1 vccd1 vccd1 _12148_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_97_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10391__C1 _10496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19744_ _19753_/CLK _19744_/D vssd1 vssd1 vccd1 vccd1 _19744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12079_ _12105_/A _12079_/B vssd1 vssd1 vccd1 vccd1 _14155_/A sky130_fd_sc_hd__nand2_2
X_16956_ _16793_/X _19386_/Q _16964_/S vssd1 vssd1 vccd1 vccd1 _16957_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10369__S0 _09632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09334__A _09819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15907_ _14847_/X _18956_/Q _15913_/S vssd1 vssd1 vccd1 vccd1 _15908_/A sky130_fd_sc_hd__mux2_1
X_19675_ _19680_/CLK _19675_/D vssd1 vssd1 vccd1 vccd1 _19675_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_38_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11486__A2 _14543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16887_ _19356_/Q _16696_/X _16891_/S vssd1 vssd1 vccd1 vccd1 _16888_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17071__A0 _16752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18626_ _19692_/CLK _18626_/D vssd1 vssd1 vccd1 vccd1 _18626_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__17610__A2 _17609_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15838_ _15838_/A vssd1 vssd1 vccd1 vccd1 _18925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18557_ _19733_/CLK _18557_/D vssd1 vssd1 vccd1 vccd1 _18557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12695__A _17882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15769_ _14879_/X _18895_/Q _15769_/S vssd1 vssd1 vccd1 vccd1 _15770_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17508_ _17508_/A vssd1 vssd1 vccd1 vccd1 _19616_/D sky130_fd_sc_hd__clkbuf_1
X_09290_ _15339_/A _11665_/B _18578_/Q vssd1 vssd1 vccd1 vccd1 _09303_/A sky130_fd_sc_hd__a21o_1
X_18488_ _19079_/CLK _18488_/D vssd1 vssd1 vccd1 vccd1 _18488_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17439_ _17439_/A vssd1 vssd1 vccd1 vccd1 _19585_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13935__A1 _10810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19109_ _19722_/CLK _19109_/D vssd1 vssd1 vccd1 vccd1 _19109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_opt_2_0_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput110 _13570_/A vssd1 vssd1 vccd1 vccd1 io_dbus_st_type[1] sky130_fd_sc_hd__buf_2
XFILLER_161_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput121 _12488_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[19] sky130_fd_sc_hd__buf_2
Xoutput132 _12503_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[29] sky130_fd_sc_hd__buf_2
Xoutput143 _11557_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wr_en sky130_fd_sc_hd__buf_2
Xoutput154 _17893_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[19] sky130_fd_sc_hd__buf_2
XFILLER_82_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput165 _17909_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[29] sky130_fd_sc_hd__buf_2
XFILLER_142_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11174__B2 _18454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10382__C1 _09247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13320__C1 _13317_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09244__A _09244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11493__B _11514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09626_ _18455_/Q vssd1 vssd1 vccd1 vccd1 _09626_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15612__A1 _15516_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09557_ _09640_/A vssd1 vssd1 vccd1 vccd1 _09649_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09898__B _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16077__A _16787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09488_ _10724_/A vssd1 vssd1 vccd1 vccd1 _10770_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_24_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10988__A1 _09177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17400__S _17402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11450_ _11434_/Y _13108_/B _11443_/X _11720_/B vssd1 vssd1 vccd1 vccd1 _11463_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10401_ _10401_/A vssd1 vssd1 vccd1 vccd1 _11112_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_20_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11381_ _18419_/Q _12555_/B _11381_/C vssd1 vssd1 vccd1 vccd1 _11381_/X sky130_fd_sc_hd__or3_1
XANTENNA__16016__S _16016_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10853__A _10950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13120_ _13365_/A vssd1 vssd1 vccd1 vccd1 _13183_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10332_ _19258_/Q _19029_/Q _18960_/Q _19354_/Q _10328_/S _09735_/A vssd1 vssd1 vccd1
+ vccd1 _10332_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09419__A _09814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13051_ _18328_/Q vssd1 vssd1 vccd1 vccd1 _13055_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15855__S _15863_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10263_ _09712_/A _10260_/X _10262_/X _09708_/X vssd1 vssd1 vccd1 vccd1 _10263_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_106_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12002_ _12186_/A vssd1 vssd1 vccd1 vccd1 _12002_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input47_A io_ibus_inst[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10194_ _18444_/Q _09309_/A _09430_/X _10193_/X vssd1 vssd1 vccd1 vccd1 _12487_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_120_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16810_ _16826_/A vssd1 vssd1 vccd1 vccd1 _16823_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__15156__A _15239_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17790_ _15146_/X _19698_/Q _17794_/S vssd1 vssd1 vccd1 vccd1 _17791_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16741_ _19306_/Q _16740_/X _16741_/S vssd1 vssd1 vccd1 vccd1 _16742_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13953_ _13952_/X _13853_/X _13995_/S vssd1 vssd1 vccd1 vccd1 _13953_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_163_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19537_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__14995__A _16718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15590__S _15590_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12904_ _12904_/A _12904_/B _12907_/B vssd1 vssd1 vccd1 vccd1 _18280_/D sky130_fd_sc_hd__nor3_1
X_19460_ _19622_/CLK _19460_/D vssd1 vssd1 vccd1 vccd1 _19460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16672_ _16672_/A vssd1 vssd1 vccd1 vccd1 _19284_/D sky130_fd_sc_hd__clkbuf_1
X_13884_ _13767_/X _13772_/X _13888_/S vssd1 vssd1 vccd1 vccd1 _13884_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15603__A1 _15503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18411_ _19788_/CLK _18411_/D vssd1 vssd1 vccd1 vccd1 _18411_/Q sky130_fd_sc_hd__dfxtp_1
X_15623_ _18830_/Q _15532_/X _15625_/S vssd1 vssd1 vccd1 vccd1 _15624_/A sky130_fd_sc_hd__mux2_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _18260_/Q _12831_/C _12834_/Y vssd1 vssd1 vccd1 vccd1 _18260_/D sky130_fd_sc_hd__o21a_1
XANTENNA__12417__A1 _19757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19391_ _19553_/CLK _19391_/D vssd1 vssd1 vccd1 vccd1 _19391_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10691__A3 _10690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _18401_/CLK _18342_/D vssd1 vssd1 vccd1 vccd1 _18342_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_178_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19442_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _16809_/A vssd1 vssd1 vccd1 vccd1 _15554_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _12766_/A vssd1 vssd1 vccd1 vccd1 _13324_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14505_ _11297_/C _18522_/Q _14565_/A vssd1 vssd1 vccd1 vccd1 _14506_/B sky130_fd_sc_hd__mux2_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _18386_/CLK _18273_/D vssd1 vssd1 vccd1 vccd1 _18273_/Q sky130_fd_sc_hd__dfxtp_1
X_11717_ _11822_/B _11715_/Y _11822_/D _11720_/B vssd1 vssd1 vccd1 vccd1 _11717_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA_clkbuf_leaf_182_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _12715_/A vssd1 vssd1 vccd1 vccd1 _18205_/A sky130_fd_sc_hd__buf_2
X_15485_ _18784_/Q _15238_/X _15485_/S vssd1 vssd1 vccd1 vccd1 _15486_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16715__A _16715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17224_ _17224_/A vssd1 vssd1 vccd1 vccd1 _19493_/D sky130_fd_sc_hd__clkbuf_1
X_11648_ _11648_/A _13650_/A vssd1 vssd1 vccd1 vccd1 _11652_/A sky130_fd_sc_hd__xnor2_1
X_14436_ _14436_/A vssd1 vssd1 vccd1 vccd1 _18490_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_101_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _18357_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput12 io_dbus_rdata[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_2
Xinput23 io_dbus_rdata[2] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_2
Xinput34 io_ibus_inst[0] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_1
X_17155_ _19473_/Q _17154_/X _17155_/S vssd1 vssd1 vccd1 vccd1 _17156_/A sky130_fd_sc_hd__mux2_1
Xinput45 io_ibus_inst[1] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10826__S1 _10740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14367_ _14366_/X _18499_/Q _14367_/S vssd1 vssd1 vccd1 vccd1 _14368_/A sky130_fd_sc_hd__mux2_1
X_11579_ _13520_/A _11599_/C _13573_/B vssd1 vssd1 vccd1 vccd1 _11579_/Y sky130_fd_sc_hd__nand3_1
Xinput56 io_ibus_inst[2] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput67 io_irq_m1_irq vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16106_ _16816_/A vssd1 vssd1 vccd1 vccd1 _16106_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13318_ _12617_/B _13311_/X _13316_/X _13317_/X vssd1 vssd1 vccd1 vccd1 _18368_/D
+ sky130_fd_sc_hd__o211a_1
X_17086_ _16774_/X _19444_/Q _17086_/S vssd1 vssd1 vccd1 vccd1 _17087_/A sky130_fd_sc_hd__mux2_1
X_14298_ _13978_/X _14300_/B _13979_/X _14297_/X vssd1 vssd1 vccd1 vccd1 _14298_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15765__S _15769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16037_ _16033_/X _19014_/Q _16049_/S vssd1 vssd1 vccd1 vccd1 _16038_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_116_clock clkbuf_opt_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _18585_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13249_ _18277_/Q _13270_/B vssd1 vssd1 vccd1 vccd1 _13249_/X sky130_fd_sc_hd__and2_1
XFILLER_124_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17988_ _19781_/Q _19780_/Q _17988_/C vssd1 vssd1 vccd1 vccd1 _17990_/B sky130_fd_sc_hd__and3_1
XFILLER_97_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19727_ _19727_/CLK _19727_/D vssd1 vssd1 vccd1 vccd1 _19727_/Q sky130_fd_sc_hd__dfxtp_1
X_16939_ _16939_/A vssd1 vssd1 vccd1 vccd1 _19378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19658_ _19725_/CLK _19658_/D vssd1 vssd1 vccd1 vccd1 _19658_/Q sky130_fd_sc_hd__dfxtp_1
X_09411_ _09411_/A vssd1 vssd1 vccd1 vccd1 _09412_/A sky130_fd_sc_hd__clkbuf_4
X_18609_ _19331_/CLK _18609_/D vssd1 vssd1 vccd1 vccd1 _18609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19589_ _19589_/CLK _19589_/D vssd1 vssd1 vccd1 vccd1 _19589_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10419__B1 _11099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ _09342_/A vssd1 vssd1 vccd1 vccd1 _11188_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__13081__A1 _19666_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09273_ _09273_/A vssd1 vssd1 vccd1 vccd1 _09274_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13984__A _13984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16360__A _16428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09673__S _09673_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12078__A1_N _14553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_80_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19804_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_130_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10950_ _10950_/A _10950_/B vssd1 vssd1 vccd1 vccd1 _10950_/X sky130_fd_sc_hd__or2_1
XFILLER_17_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_95_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19779_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09609_ _09734_/A vssd1 vssd1 vccd1 vccd1 _10131_/S sky130_fd_sc_hd__buf_4
XANTENNA__11951__B _13620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10881_ _12465_/A _10834_/X _12466_/A _11779_/A vssd1 vssd1 vccd1 vccd1 _10881_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15061__A2 _13422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12620_ _19811_/Q vssd1 vssd1 vccd1 vccd1 _18075_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ _19776_/Q _12548_/X _12666_/B vssd1 vssd1 vccd1 vccd1 _12551_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14754__S _14762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17130__S _17130_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11502_ _18581_/Q vssd1 vssd1 vccd1 vccd1 _14580_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_129_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15270_ _18689_/Q _15133_/X _15278_/S vssd1 vssd1 vccd1 vccd1 _15271_/A sky130_fd_sc_hd__mux2_1
X_12482_ _12482_/A _12483_/B vssd1 vssd1 vccd1 vccd1 _12482_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11433_ _12555_/B _18417_/Q _11427_/X _11432_/X vssd1 vssd1 vccd1 vccd1 _11463_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_14221_ _13909_/X _14219_/X _14220_/Y _15123_/A vssd1 vssd1 vccd1 vccd1 _14221_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_137_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11386__A1 _18427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19591_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09149__A _09149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14152_ _14297_/A _14155_/A vssd1 vssd1 vccd1 vccd1 _14152_/X sky130_fd_sc_hd__or2_1
XFILLER_153_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11364_ _11372_/A _11584_/A vssd1 vssd1 vccd1 vccd1 _13584_/C sky130_fd_sc_hd__and2_2
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17510__A1 _16705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13103_ _18345_/Q _12731_/X _13101_/X _13102_/X vssd1 vssd1 vccd1 vccd1 _18345_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10315_ _18864_/Q _19322_/Q _11157_/S vssd1 vssd1 vccd1 vccd1 _10315_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14083_ _11956_/X _14070_/X _14082_/X _13828_/X vssd1 vssd1 vccd1 vccd1 _14083_/X
+ sky130_fd_sc_hd__a211o_1
X_18960_ _19549_/CLK _18960_/D vssd1 vssd1 vccd1 vccd1 _18960_/Q sky130_fd_sc_hd__dfxtp_1
X_11295_ _14513_/A _14511_/A _11297_/B _11297_/C vssd1 vssd1 vccd1 vccd1 _11468_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17911_ _19758_/Q _12186_/A _12437_/X _12440_/X _17895_/X vssd1 vssd1 vccd1 vccd1
+ _19758_/D sky130_fd_sc_hd__o221a_1
X_13034_ _13034_/A _13034_/B _13034_/C vssd1 vssd1 vccd1 vccd1 _18323_/D sky130_fd_sc_hd__nor3_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10246_ _18770_/Q _18999_/Q _18930_/Q _19228_/Q _10279_/S _10245_/X vssd1 vssd1 vccd1
+ vccd1 _10246_/X sky130_fd_sc_hd__mux4_1
X_18891_ _19543_/CLK _18891_/D vssd1 vssd1 vccd1 vccd1 _18891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_129_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_48_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19556_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17842_ _17842_/A vssd1 vssd1 vccd1 vccd1 _19721_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10897__B1 _10774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10177_ _10177_/A _10177_/B vssd1 vssd1 vccd1 vccd1 _10177_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17773_ _17773_/A vssd1 vssd1 vccd1 vccd1 _19690_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14985_ _16715_/A vssd1 vssd1 vccd1 vccd1 _16819_/A sky130_fd_sc_hd__buf_2
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19512_ _19608_/CLK _19512_/D vssd1 vssd1 vccd1 vccd1 _19512_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09503__A1 _09486_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16724_ _16724_/A vssd1 vssd1 vccd1 vccd1 _19300_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17305__S _17313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13936_ _13939_/B _13936_/B vssd1 vssd1 vccd1 vccd1 _13943_/B sky130_fd_sc_hd__nand2_1
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12957__B _18295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19443_ _19704_/CLK _19443_/D vssd1 vssd1 vccd1 vccd1 _19443_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09612__A _10177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16655_ _19279_/Q _16654_/X _16655_/S vssd1 vssd1 vccd1 vccd1 _16656_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13867_ _13745_/X _13665_/X _14314_/A _13866_/X vssd1 vssd1 vccd1 vccd1 _13868_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15606_ _18822_/Q _15506_/X _15614_/S vssd1 vssd1 vccd1 vccd1 _15607_/A sky130_fd_sc_hd__mux2_1
X_12818_ _12821_/B _12821_/C _12817_/X vssd1 vssd1 vccd1 vccd1 _12818_/Y sky130_fd_sc_hd__a21oi_1
X_19374_ _19691_/CLK _19374_/D vssd1 vssd1 vccd1 vccd1 _19374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16586_ _16586_/A vssd1 vssd1 vccd1 vccd1 _19248_/D sky130_fd_sc_hd__clkbuf_1
X_13798_ _14089_/A vssd1 vssd1 vccd1 vccd1 _14212_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18325_ _18330_/CLK _18325_/D vssd1 vssd1 vccd1 vccd1 _18325_/Q sky130_fd_sc_hd__dfxtp_1
X_15537_ _15537_/A vssd1 vssd1 vccd1 vccd1 _18799_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _12749_/A vssd1 vssd1 vccd1 vccd1 _12749_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12973__A _12983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18256_ _19855_/CLK _18256_/D vssd1 vssd1 vccd1 vccd1 _18256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15468_ _18776_/Q _15213_/X _15470_/S vssd1 vssd1 vccd1 vccd1 _15469_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17207_ _17207_/A vssd1 vssd1 vccd1 vccd1 _19488_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11589__A _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14563__A1 _18574_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14419_ _15027_/A _18517_/Q _14424_/S vssd1 vssd1 vccd1 vccd1 _14420_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18187_ _19849_/Q _18185_/B _18186_/Y vssd1 vssd1 vccd1 vccd1 _19849_/D sky130_fd_sc_hd__o21a_1
XFILLER_129_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15399_ _15399_/A vssd1 vssd1 vccd1 vccd1 _18746_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09665__S1 _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17138_ _13203_/X _15241_/X _17137_/X _15243_/Y vssd1 vssd1 vccd1 vccd1 _17226_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_116_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09960_ _09969_/A _09960_/B vssd1 vssd1 vccd1 vccd1 _09960_/X sky130_fd_sc_hd__or2_1
X_17069_ _16749_/X _19436_/Q _17075_/S vssd1 vssd1 vccd1 vccd1 _17070_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09891_ _19654_/Q _19071_/Q _19108_/Q _18714_/Q _09809_/X _09881_/X vssd1 vssd1 vccd1
+ vccd1 _09891_/X sky130_fd_sc_hd__mux4_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12213__A _14211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17568__A1 _16790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09522__A _09522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10668__A _10668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09325_ _10640_/A vssd1 vssd1 vccd1 vccd1 _10524_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09256_ _16212_/B _11519_/A _18569_/Q vssd1 vssd1 vccd1 vccd1 _11368_/A sky130_fd_sc_hd__a21o_1
XFILLER_167_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13698__B _13720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09187_ _10107_/A vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10040__A1 _09892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14306__A1 _14305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10100_ _10100_/A vssd1 vssd1 vccd1 vccd1 _10102_/A sky130_fd_sc_hd__inv_2
XFILLER_89_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11080_ _10601_/X _11080_/B _11080_/C vssd1 vssd1 vccd1 vccd1 _11244_/B sky130_fd_sc_hd__and3b_1
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_130_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14322__B _14324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ _18870_/Q _19328_/Q _10033_/S vssd1 vssd1 vccd1 vccd1 _10032_/B sky130_fd_sc_hd__mux2_1
XFILLER_103_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10974__S0 _10668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14770_ input28/X _14703_/A _14769_/X _14732_/X vssd1 vssd1 vccd1 vccd1 _16657_/A
+ sky130_fd_sc_hd__a22o_1
X_11982_ _19740_/Q vssd1 vssd1 vccd1 vccd1 _17878_/A sky130_fd_sc_hd__buf_4
XFILLER_57_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13721_ _14003_/A vssd1 vssd1 vccd1 vccd1 _13721_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10933_ _09481_/A _10933_/B vssd1 vssd1 vccd1 vccd1 _10933_/X sky130_fd_sc_hd__and2b_1
XANTENNA__16964__S _16964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16440_ _16045_/X _19182_/Q _16442_/S vssd1 vssd1 vccd1 vccd1 _16441_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13652_ _13641_/X _13649_/X _13968_/S vssd1 vssd1 vccd1 vccd1 _13652_/X sky130_fd_sc_hd__mux2_1
X_10864_ _10859_/X _10861_/Y _09224_/A _10863_/Y vssd1 vssd1 vccd1 vccd1 _10864_/X
+ sky130_fd_sc_hd__a211o_1
X_12603_ _12603_/A vssd1 vssd1 vccd1 vccd1 _12604_/A sky130_fd_sc_hd__clkbuf_2
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _16428_/S vssd1 vssd1 vccd1 vccd1 _16380_/S sky130_fd_sc_hd__buf_2
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10795_ _10844_/A _10795_/B vssd1 vssd1 vccd1 vccd1 _10795_/X sky130_fd_sc_hd__or2_1
X_13583_ _13583_/A _13583_/B vssd1 vssd1 vccd1 vccd1 _13585_/C sky130_fd_sc_hd__nor2_1
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18110_ _19824_/Q _18110_/B _18110_/C vssd1 vssd1 vccd1 vccd1 _18111_/C sky130_fd_sc_hd__and3_1
XFILLER_9_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15322_ _18713_/Q _15216_/X _15322_/S vssd1 vssd1 vccd1 vccd1 _15323_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_55_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12534_ _12545_/A vssd1 vssd1 vccd1 vccd1 _12566_/A sky130_fd_sc_hd__inv_2
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19090_ _19635_/CLK _19090_/D vssd1 vssd1 vccd1 vccd1 _19090_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13348__A2 _13346_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18041_ _18043_/A _18043_/C _18040_/Y vssd1 vssd1 vccd1 vccd1 _19799_/D sky130_fd_sc_hd__o21a_1
X_15253_ _15253_/A vssd1 vssd1 vccd1 vccd1 _18685_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12465_ _12465_/A _12469_/B vssd1 vssd1 vccd1 vccd1 _12465_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14204_ _13943_/A _14199_/Y _14203_/Y vssd1 vssd1 vccd1 vccd1 _14204_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11202__A _11202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11416_ _18543_/Q vssd1 vssd1 vccd1 vccd1 _12540_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15184_ _16686_/A vssd1 vssd1 vccd1 vccd1 _15184_/X sky130_fd_sc_hd__clkbuf_2
X_12396_ _14584_/A _13525_/A _12345_/X _12503_/A vssd1 vssd1 vccd1 vccd1 _12397_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_153_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14135_ _14135_/A _14135_/B vssd1 vssd1 vccd1 vccd1 _14135_/Y sky130_fd_sc_hd__nand2_1
X_11347_ _11358_/B _11642_/C vssd1 vssd1 vccd1 vccd1 _11347_/Y sky130_fd_sc_hd__nor2_2
XFILLER_126_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14066_ _13949_/A _14063_/X _14065_/Y _13950_/X vssd1 vssd1 vccd1 vccd1 _14066_/X
+ sky130_fd_sc_hd__a211o_1
X_18943_ _19337_/CLK _18943_/D vssd1 vssd1 vccd1 vccd1 _18943_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output78_A _12041_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ _11220_/Y _11249_/A _11223_/X _11224_/Y _11277_/X vssd1 vssd1 vccd1 vccd1
+ _11278_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_79_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13017_ _18316_/Q _18318_/Q _18317_/Q _13017_/D vssd1 vssd1 vccd1 vccd1 _13026_/D
+ sky130_fd_sc_hd__and4_1
X_10229_ _11119_/A _10229_/B vssd1 vssd1 vccd1 vccd1 _10229_/Y sky130_fd_sc_hd__nor2_1
X_18874_ _19556_/CLK _18874_/D vssd1 vssd1 vccd1 vccd1 _18874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11575__C _15095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17825_ _15197_/X _19714_/Q _17827_/S vssd1 vssd1 vccd1 vccd1 _17826_/A sky130_fd_sc_hd__mux2_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17756_ _18486_/Q _17757_/B vssd1 vssd1 vccd1 vccd1 _17765_/C sky130_fd_sc_hd__or2_1
X_14968_ _17728_/A _14979_/C vssd1 vssd1 vccd1 vccd1 _14978_/B sky130_fd_sc_hd__and2_1
X_16707_ _19295_/Q _16705_/X _16719_/S vssd1 vssd1 vccd1 vccd1 _16708_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09342__A _09342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10098__B2 _18446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13919_ _14135_/A _13889_/X _13816_/X vssd1 vssd1 vccd1 vccd1 _13919_/X sky130_fd_sc_hd__o21a_1
X_17687_ _17707_/A vssd1 vssd1 vccd1 vccd1 _17718_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__16874__S _16880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14899_ _14838_/X _14897_/X _14898_/X vssd1 vssd1 vccd1 vccd1 _14899_/Y sky130_fd_sc_hd__a21oi_1
X_19426_ _19720_/CLK _19426_/D vssd1 vssd1 vccd1 vccd1 _19426_/Q sky130_fd_sc_hd__dfxtp_1
X_16638_ _16638_/A vssd1 vssd1 vccd1 vccd1 _19274_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15981__A0 _14808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19357_ _19616_/CLK _19357_/D vssd1 vssd1 vccd1 vccd1 _19357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16569_ _19240_/Q _15583_/X _16569_/S vssd1 vssd1 vccd1 vccd1 _16570_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09110_ _11317_/A vssd1 vssd1 vccd1 vccd1 _11472_/A sky130_fd_sc_hd__buf_2
XFILLER_148_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18308_ _18329_/CLK _18308_/D vssd1 vssd1 vccd1 vccd1 _18308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19288_ _19709_/CLK _19288_/D vssd1 vssd1 vccd1 vccd1 _19288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18239_ _19868_/Q _18239_/B _18239_/C vssd1 vssd1 vccd1 vccd1 _18241_/B sky130_fd_sc_hd__and3_1
XANTENNA__14536__A1 _16919_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09963__A1 _09892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09943_ _19652_/Q _19069_/Q _19106_/Q _18712_/Q _09866_/X _09869_/X vssd1 vssd1 vccd1
+ vccd1 _09944_/B sky130_fd_sc_hd__mux4_2
XANTENNA__11766__B _15255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17238__A0 _18455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09874_ _18611_/Q _19300_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09875_/B sky130_fd_sc_hd__mux2_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14674__A1_N input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13473__S _13475_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15254__A _17762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09877__S1 _09810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09308_ _09308_/A vssd1 vssd1 vccd1 vccd1 _09309_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_139_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10580_ _09515_/A _10580_/B vssd1 vssd1 vccd1 vccd1 _10580_/X sky130_fd_sc_hd__and2b_1
XFILLER_142_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_7_0_clock clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_139_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14527__A1 _11511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09239_ _19628_/Q _19466_/Q _18912_/Q _18682_/Q _09190_/A _09149_/A vssd1 vssd1 vccd1
+ vccd1 _09240_/B sky130_fd_sc_hd__mux4_1
XFILLER_10_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12118__A _19745_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11022__A _18427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12250_ _18372_/Q _12272_/C vssd1 vssd1 vccd1 vccd1 _12250_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10013__A1 _09783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11201_ _09901_/Y _11152_/Y _11198_/Y _11199_/Y _11251_/A vssd1 vssd1 vccd1 vccd1
+ _11220_/B sky130_fd_sc_hd__a311o_1
XANTENNA__11957__A _19739_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12181_ _12181_/A _14203_/B vssd1 vssd1 vccd1 vccd1 _12182_/B sky130_fd_sc_hd__nor2_1
XFILLER_163_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11761__A1 _18415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11132_ _11132_/A vssd1 vssd1 vccd1 vccd1 _11132_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17229__A0 _18452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15863__S _15863_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15940_ _15022_/X _18971_/Q _15946_/S vssd1 vssd1 vccd1 vccd1 _15941_/A sky130_fd_sc_hd__mux2_1
X_11063_ _19597_/Q _19435_/Q _18881_/Q _18651_/Q _10932_/S _10772_/A vssd1 vssd1 vccd1
+ vccd1 _11063_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10947__S0 _10719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10014_ _19424_/Q _19200_/Q _19717_/Q _19168_/Q _09782_/A _09979_/X vssd1 vssd1 vccd1
+ vccd1 _10014_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15871_ _15871_/A vssd1 vssd1 vccd1 vccd1 _18940_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17610_ _15258_/X _17609_/Y _15255_/B vssd1 vssd1 vccd1 vccd1 _17610_/X sky130_fd_sc_hd__a21o_1
XFILLER_64_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14822_ _14821_/X _18595_/Q _14822_/S vssd1 vssd1 vccd1 vccd1 _14823_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13266__A1 _12727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18590_ _19698_/CLK _18590_/D vssd1 vssd1 vccd1 vccd1 _18590_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14463__A0 _18503_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17541_ _17541_/A vssd1 vssd1 vccd1 vccd1 _19630_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09565__S0 _09553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14753_ _16755_/A vssd1 vssd1 vccd1 vccd1 _14753_/X sky130_fd_sc_hd__clkbuf_2
X_11965_ _19739_/Q _11928_/X _11960_/X _11964_/X vssd1 vssd1 vccd1 vccd1 _17876_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__16694__S _16703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13704_ _13891_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13706_/A sky130_fd_sc_hd__and2_1
X_17472_ _19600_/Q _16651_/X _17474_/S vssd1 vssd1 vccd1 vccd1 _17473_/A sky130_fd_sc_hd__mux2_1
X_10916_ _10956_/A _10913_/X _10915_/X _09223_/A vssd1 vssd1 vccd1 vccd1 _10917_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14684_ _14580_/A _14633_/X _14680_/X input53/X vssd1 vssd1 vccd1 vccd1 _14685_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11896_ _10601_/B _18499_/Q _11948_/A vssd1 vssd1 vccd1 vccd1 _13614_/A sky130_fd_sc_hd__mux2_8
XFILLER_72_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19211_ _19696_/CLK _19211_/D vssd1 vssd1 vccd1 vccd1 _19211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16423_ _16423_/A vssd1 vssd1 vccd1 vccd1 _19175_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11029__B1 _09177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13635_ _13631_/X _13633_/X _13741_/S vssd1 vssd1 vccd1 vccd1 _13635_/X sky130_fd_sc_hd__mux2_1
X_10847_ _19634_/Q _19051_/Q _19088_/Q _18694_/Q _10648_/S _10634_/A vssd1 vssd1 vccd1
+ vccd1 _10848_/B sky130_fd_sc_hd__mux4_1
XANTENNA__11124__S0 _10279_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19142_ _19723_/CLK _19142_/D vssd1 vssd1 vccd1 vccd1 _19142_/Q sky130_fd_sc_hd__dfxtp_1
X_16354_ _16354_/A vssd1 vssd1 vccd1 vccd1 _19145_/D sky130_fd_sc_hd__clkbuf_1
X_13566_ _15116_/A vssd1 vssd1 vccd1 vccd1 _13566_/X sky130_fd_sc_hd__buf_2
XFILLER_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10778_ _10807_/A _10778_/B vssd1 vssd1 vccd1 vccd1 _10778_/X sky130_fd_sc_hd__or2_1
XFILLER_40_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15305_ _18705_/Q _15191_/X _15311_/S vssd1 vssd1 vccd1 vccd1 _15306_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12517_ _12664_/A vssd1 vssd1 vccd1 vccd1 _12518_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10252__B2 _10251_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19073_ _19723_/CLK _19073_/D vssd1 vssd1 vccd1 vccd1 _19073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16285_ _17391_/B _17064_/B vssd1 vssd1 vccd1 vccd1 _16342_/A sky130_fd_sc_hd__or2_2
X_13497_ _18407_/Q _12779_/X _13497_/S vssd1 vssd1 vccd1 vccd1 _13498_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18024_ _18023_/A _18023_/B _19794_/Q vssd1 vssd1 vccd1 vccd1 _18025_/C sky130_fd_sc_hd__a21oi_1
XFILLER_117_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15236_ _18681_/Q _15235_/X _15239_/S vssd1 vssd1 vccd1 vccd1 _15237_/A sky130_fd_sc_hd__mux2_1
X_12448_ _14324_/A _12422_/B _13702_/A vssd1 vssd1 vccd1 vccd1 _12449_/B sky130_fd_sc_hd__o21ai_1
XFILLER_125_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15339__A _15339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15167_ _15167_/A vssd1 vssd1 vccd1 vccd1 _18659_/D sky130_fd_sc_hd__clkbuf_1
X_12379_ _14300_/A _12379_/B vssd1 vssd1 vccd1 vccd1 _12383_/A sky130_fd_sc_hd__xnor2_1
XFILLER_5_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09337__A _10706_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14118_ _18439_/Q _14117_/X _14209_/S vssd1 vssd1 vccd1 vccd1 _14119_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15098_ _18624_/Q _13566_/X _15097_/X _11779_/Y vssd1 vssd1 vccd1 vccd1 _18624_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16869__S _16869_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18926_ _19640_/CLK _18926_/D vssd1 vssd1 vccd1 vccd1 _18926_/Q sky130_fd_sc_hd__dfxtp_1
X_14049_ _13726_/X _14036_/X _14048_/X _14012_/X vssd1 vssd1 vccd1 vccd1 _14049_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_122_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09771__S _10010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10938__S0 _10706_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18857_ _19541_/CLK _18857_/D vssd1 vssd1 vccd1 vccd1 _18857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09590_ _09728_/A vssd1 vssd1 vccd1 vccd1 _09595_/A sky130_fd_sc_hd__clkbuf_4
X_17808_ _15171_/X _19706_/Q _17816_/S vssd1 vssd1 vccd1 vccd1 _17809_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13257__A1 _19834_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18788_ _19691_/CLK _18788_/D vssd1 vssd1 vccd1 vccd1 _18788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17739_ _17743_/B _17738_/Y _17711_/X vssd1 vssd1 vccd1 vccd1 _17739_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09556__S0 _09553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11807__A2 _11740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10166__S1 _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11107__A _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19409_ _19571_/CLK _19409_/D vssd1 vssd1 vccd1 vccd1 _19409_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14757__A1 _13181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15948__S _15950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15182__A1 _15181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09247__A _09247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16779__S _16791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09926_ _09926_/A vssd1 vssd1 vccd1 vccd1 _09927_/A sky130_fd_sc_hd__buf_2
XANTENNA__17464__A _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09857_ _19654_/Q _19071_/Q _19108_/Q _18714_/Q _09163_/A _09843_/A vssd1 vssd1 vccd1
+ vccd1 _09858_/B sky130_fd_sc_hd__mux4_1
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _09788_/A _09788_/B vssd1 vssd1 vccd1 vccd1 _09788_/X sky130_fd_sc_hd__or2_1
XFILLER_46_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12401__A _12401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _12016_/S vssd1 vssd1 vccd1 vccd1 _12119_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10482__A1 _09212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10701_ _10701_/A _10701_/B vssd1 vssd1 vccd1 vccd1 _10701_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10880__A1_N _18431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11994_/A vssd1 vssd1 vccd1 vccd1 _17241_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__16019__S _16027_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11106__S0 _10230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13420_ _18265_/Q _12582_/X _12584_/X _19854_/Q _13419_/X vssd1 vssd1 vccd1 vccd1
+ _13420_/X sky130_fd_sc_hd__a221o_1
XANTENNA__13232__A _17781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10632_ _10712_/A vssd1 vssd1 vccd1 vccd1 _10785_/A sky130_fd_sc_hd__buf_2
XFILLER_139_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17698__A0 _12598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10234__A1 _10219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13351_ _12757_/X _13139_/X _13349_/X _13350_/X vssd1 vssd1 vccd1 vccd1 _18373_/D
+ sky130_fd_sc_hd__o211a_1
X_10563_ _10559_/X _10561_/X _10562_/X _10574_/A _09434_/A vssd1 vssd1 vccd1 vccd1
+ _10568_/B sky130_fd_sc_hd__o221a_1
XFILLER_155_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14762__S _14762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12302_ _14575_/A _12344_/A _12345_/A _12499_/A vssd1 vssd1 vccd1 vccd1 _12303_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_16070_ _16070_/A vssd1 vssd1 vccd1 vccd1 _19024_/D sky130_fd_sc_hd__clkbuf_1
X_13282_ _14514_/A vssd1 vssd1 vccd1 vccd1 _13282_/X sky130_fd_sc_hd__buf_2
XFILLER_6_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10494_ _10494_/A _10494_/B _10494_/C vssd1 vssd1 vccd1 vccd1 _10494_/X sky130_fd_sc_hd__or3_4
XANTENNA__12790__B _16847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15021_ _16725_/A vssd1 vssd1 vccd1 vccd1 _16829_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15159__A _16661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12233_ _12233_/A _13615_/A vssd1 vssd1 vccd1 vccd1 _12234_/A sky130_fd_sc_hd__xnor2_1
XFILLER_108_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11195__C1 _09394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12164_ _19747_/Q _12215_/C vssd1 vssd1 vccd1 vccd1 _12164_/X sky130_fd_sc_hd__xor2_1
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11115_ _10392_/A _11114_/X _09529_/X vssd1 vssd1 vccd1 vccd1 _11115_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_151_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16972_ _16972_/A vssd1 vssd1 vccd1 vccd1 _19393_/D sky130_fd_sc_hd__clkbuf_1
X_19760_ _19866_/CLK _19760_/D vssd1 vssd1 vccd1 vccd1 _19760_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_150_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12095_ _12095_/A _12095_/B _12117_/C vssd1 vssd1 vccd1 vccd1 _12095_/Y sky130_fd_sc_hd__nand3_1
XFILLER_150_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18711_ _19718_/CLK _18711_/D vssd1 vssd1 vccd1 vccd1 _18711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11046_ _11046_/A _11046_/B vssd1 vssd1 vccd1 vccd1 _11046_/Y sky130_fd_sc_hd__nand2_1
X_15923_ _15923_/A vssd1 vssd1 vccd1 vccd1 _18963_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19691_ _19691_/CLK _19691_/D vssd1 vssd1 vccd1 vccd1 _19691_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10396__S1 _09602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18642_ _19628_/CLK _18642_/D vssd1 vssd1 vccd1 vccd1 _18642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13239__A1 _19668_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15854_ _15865_/A vssd1 vssd1 vccd1 vccd1 _15863_/S sky130_fd_sc_hd__buf_4
XFILLER_37_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14805_ input31/X _14801_/X _14804_/X vssd1 vssd1 vccd1 vccd1 _14805_/X sky130_fd_sc_hd__a21o_1
XFILLER_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18573_ _18578_/CLK _18573_/D vssd1 vssd1 vccd1 vccd1 _18573_/Q sky130_fd_sc_hd__dfxtp_1
X_15785_ _14964_/X _18902_/Q _15791_/S vssd1 vssd1 vccd1 vccd1 _15786_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12997_ _12997_/A _13003_/C vssd1 vssd1 vccd1 vccd1 _12997_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__16718__A _16718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17524_ _17524_/A vssd1 vssd1 vccd1 vccd1 _19623_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17313__S _17313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14736_ _15018_/A _13163_/B _14735_/X vssd1 vssd1 vccd1 vccd1 _14736_/X sky130_fd_sc_hd__a21o_2
X_11948_ _11948_/A vssd1 vssd1 vccd1 vccd1 _12060_/A sky130_fd_sc_hd__buf_2
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10473__A1 _09212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ _16835_/X _19593_/Q _17457_/S vssd1 vssd1 vccd1 vccd1 _17456_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14667_ _14667_/A vssd1 vssd1 vccd1 vccd1 _18575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11879_ _11879_/A _11879_/B vssd1 vssd1 vccd1 vccd1 _11880_/A sky130_fd_sc_hd__xnor2_4
XFILLER_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16406_ _16406_/A vssd1 vssd1 vccd1 vccd1 _19167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13618_ _14026_/B _12262_/B _13685_/S vssd1 vssd1 vccd1 vccd1 _13618_/X sky130_fd_sc_hd__mux2_1
X_17386_ _17386_/A vssd1 vssd1 vccd1 vccd1 _19562_/D sky130_fd_sc_hd__clkbuf_1
X_14598_ input45/X vssd1 vssd1 vccd1 vccd1 _14598_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19125_ _19639_/CLK _19125_/D vssd1 vssd1 vccd1 vccd1 _19125_/Q sky130_fd_sc_hd__dfxtp_1
X_16337_ _16337_/A vssd1 vssd1 vccd1 vccd1 _19137_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13549_ _13549_/A vssd1 vssd1 vccd1 vccd1 _18420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09766__S _10010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19056_ _19706_/CLK _19056_/D vssd1 vssd1 vccd1 vccd1 _19056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16268_ _16112_/X _19107_/Q _16268_/S vssd1 vssd1 vccd1 vccd1 _16269_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18007_ _18033_/A _18007_/B _18011_/C vssd1 vssd1 vccd1 vccd1 _19787_/D sky130_fd_sc_hd__nor3_1
XFILLER_133_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15219_ _16721_/A vssd1 vssd1 vccd1 vccd1 _15219_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15069__A _18489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14911__A1 _12594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16199_ _16119_/X _19072_/Q _16205_/S vssd1 vssd1 vccd1 vccd1 _16200_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10528__A2 _10518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13478__A1 _13307_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_177_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ _19655_/Q _19072_/Q _19109_/Q _18715_/Q _10257_/S _10080_/A vssd1 vssd1 vccd1
+ vccd1 _09712_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09777__S0 _09760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18909_ _19271_/CLK _18909_/D vssd1 vssd1 vccd1 vccd1 _18909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09642_ _09642_/A _09642_/B vssd1 vssd1 vccd1 vccd1 _09642_/X sky130_fd_sc_hd__and2_1
XFILLER_82_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14427__A0 _18488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09573_ _09214_/A _09566_/X _09568_/X _09572_/X _09247_/A vssd1 vssd1 vccd1 vccd1
+ _09573_/X sky130_fd_sc_hd__a311o_4
XANTENNA__10139__S1 _09867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12989__B1 _12922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15532__A _16787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10216__A1 _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13469__A1 _12713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09909_ _09919_/A _09906_/X _09908_/X _09231_/A vssd1 vssd1 vccd1 vccd1 _09909_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10378__S1 _10349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12920_ _12943_/A _12920_/B _12930_/D vssd1 vssd1 vccd1 vccd1 _18284_/D sky130_fd_sc_hd__nor3_1
XANTENNA__10350__S _10350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12851_ _12851_/A _12851_/B _12851_/C vssd1 vssd1 vccd1 vccd1 _18265_/D sky130_fd_sc_hd__nor3_1
XFILLER_132_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11970__A _11970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11802_ _11790_/X _11796_/X _11800_/X _11801_/X vssd1 vssd1 vccd1 vccd1 _11803_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15570_ _16825_/A vssd1 vssd1 vccd1 vccd1 _15570_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _12731_/X _12765_/X _12781_/X _12763_/X vssd1 vssd1 vccd1 vccd1 _18300_/D
+ sky130_fd_sc_hd__o22a_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _14577_/A vssd1 vssd1 vccd1 vccd1 _14572_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10455__A1 _10395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _11776_/A _11733_/B vssd1 vssd1 vccd1 vccd1 _11741_/A sky130_fd_sc_hd__nor2_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _17240_/A vssd1 vssd1 vccd1 vccd1 _19498_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _18498_/Q _11901_/A _14454_/S vssd1 vssd1 vccd1 vccd1 _14453_/A sky130_fd_sc_hd__mux2_1
X_11664_ _11664_/A _11664_/B _11664_/C _11664_/D vssd1 vssd1 vccd1 vccd1 _11665_/D
+ sky130_fd_sc_hd__or4_1
XANTENNA__10207__A1 _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13403_ _13403_/A hold3/A vssd1 vssd1 vccd1 vccd1 _13403_/Y sky130_fd_sc_hd__nand2_1
XFILLER_168_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17171_ _18435_/Q _13245_/X _17184_/S vssd1 vssd1 vccd1 vccd1 _17171_/X sky130_fd_sc_hd__mux2_1
X_10615_ _10960_/A vssd1 vssd1 vccd1 vccd1 _10906_/A sky130_fd_sc_hd__clkbuf_4
X_14383_ _18473_/Q vssd1 vssd1 vccd1 vccd1 _14883_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11595_ _11591_/Y _18490_/Q _11697_/S vssd1 vssd1 vccd1 vccd1 _12510_/B sky130_fd_sc_hd__mux2_8
XANTENNA__10758__A2 _10748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16122_ _16832_/A vssd1 vssd1 vccd1 vccd1 _16122_/X sky130_fd_sc_hd__clkbuf_1
X_13334_ _13297_/X _13325_/Y _13333_/X _13306_/X _18640_/Q vssd1 vssd1 vccd1 vccd1
+ _13334_/X sky130_fd_sc_hd__a32o_4
X_10546_ _10739_/A vssd1 vssd1 vccd1 vccd1 _10813_/A sky130_fd_sc_hd__buf_2
Xclkbuf_3_4_0_clock clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_109_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16894__A1 _16705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16053_ _16051_/X _19019_/Q _16065_/S vssd1 vssd1 vccd1 vccd1 _16054_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13265_ _13265_/A _13295_/B vssd1 vssd1 vccd1 vccd1 _13265_/X sky130_fd_sc_hd__or2_1
XFILLER_157_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10477_ _10477_/A _10477_/B vssd1 vssd1 vccd1 vccd1 _10477_/X sky130_fd_sc_hd__or2_1
XFILLER_136_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15004_ _15015_/B _15003_/Y _14737_/A vssd1 vssd1 vccd1 vccd1 _15004_/Y sky130_fd_sc_hd__o21ai_1
X_12216_ _19749_/Q _12217_/B vssd1 vssd1 vccd1 vccd1 _12218_/A sky130_fd_sc_hd__nor2_1
XFILLER_155_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13196_ _18624_/Q _13196_/B vssd1 vssd1 vccd1 vccd1 _13196_/X sky130_fd_sc_hd__or2_1
XFILLER_123_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12380__A1 _18518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19812_ _19812_/CLK _19812_/D vssd1 vssd1 vccd1 vccd1 _19812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12147_ _19677_/Q _12191_/A _17221_/A vssd1 vssd1 vccd1 vccd1 _12147_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10554__A_N _12476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19743_ _19753_/CLK _19743_/D vssd1 vssd1 vccd1 vccd1 _19743_/Q sky130_fd_sc_hd__dfxtp_4
X_16955_ _16977_/A vssd1 vssd1 vccd1 vccd1 _16964_/S sky130_fd_sc_hd__buf_4
X_12078_ _14553_/A _12026_/A _12005_/A _12485_/A vssd1 vssd1 vccd1 vccd1 _12079_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15906_ _15906_/A vssd1 vssd1 vccd1 vccd1 _18955_/D sky130_fd_sc_hd__clkbuf_1
X_11029_ _09169_/A _11028_/X _09177_/A vssd1 vssd1 vccd1 vccd1 _11029_/X sky130_fd_sc_hd__a21o_1
X_19674_ _19682_/CLK _19674_/D vssd1 vssd1 vccd1 vccd1 _19674_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__12041__A _12041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16886_ _16886_/A vssd1 vssd1 vccd1 vccd1 _19355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15837_ _14856_/X _18925_/Q _15841_/S vssd1 vssd1 vccd1 vccd1 _15838_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18625_ _19692_/CLK _18625_/D vssd1 vssd1 vccd1 vccd1 _18625_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__11891__B1 _11901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12976__A _12997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17043__S _17047_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11880__A _11880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18556_ _19733_/CLK _18556_/D vssd1 vssd1 vccd1 vccd1 _18556_/Q sky130_fd_sc_hd__dfxtp_1
X_15768_ _15768_/A vssd1 vssd1 vccd1 vccd1 _18894_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14719_ _16138_/A _16138_/B _15960_/C vssd1 vssd1 vccd1 vccd1 _17391_/A sky130_fd_sc_hd__or3_4
X_17507_ _19616_/Q _16702_/X _17507_/S vssd1 vssd1 vccd1 vccd1 _17508_/A sky130_fd_sc_hd__mux2_1
X_18487_ _18487_/CLK _18487_/D vssd1 vssd1 vccd1 vccd1 _18487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15699_ _15721_/A vssd1 vssd1 vccd1 vccd1 _15708_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_21_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10496__A _10496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17438_ _16809_/X _19585_/Q _17446_/S vssd1 vssd1 vccd1 vccd1 _17439_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17369_ _17369_/A vssd1 vssd1 vccd1 vccd1 _19554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19108_ _19721_/CLK _19108_/D vssd1 vssd1 vccd1 vccd1 _19108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19039_ _19721_/CLK _19039_/D vssd1 vssd1 vccd1 vccd1 _19039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12216__A _19749_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput100 _11787_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[5] sky130_fd_sc_hd__buf_2
Xoutput111 _12459_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[0] sky130_fd_sc_hd__buf_2
Xoutput122 _12461_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[1] sky130_fd_sc_hd__buf_2
Xoutput133 _12462_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[2] sky130_fd_sc_hd__buf_2
XFILLER_161_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput144 _11572_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[0] sky130_fd_sc_hd__buf_2
Xoutput155 _17857_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[1] sky130_fd_sc_hd__buf_2
XFILLER_142_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput166 _11685_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[2] sky130_fd_sc_hd__buf_2
XANTENNA__11174__A2 _11164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14431__A _14431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09525__A _10387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09625_ _09625_/A vssd1 vssd1 vccd1 vccd1 _09625_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_16_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16358__A _16503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15262__A _15262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ _19432_/Q _19208_/Q _19725_/Q _19176_/Q _09553_/X _09555_/X vssd1 vssd1 vccd1
+ vccd1 _09556_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13084__C1 _13083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09487_ _18977_/Q vssd1 vssd1 vccd1 vccd1 _10724_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15376__A1 _15187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11014__B _11014_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15201__S _15201_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10400_ _10400_/A _10400_/B vssd1 vssd1 vccd1 vccd1 _10400_/Y sky130_fd_sc_hd__nor2_1
X_11380_ _18418_/Q vssd1 vssd1 vccd1 vccd1 _12555_/B sky130_fd_sc_hd__buf_2
XANTENNA__15128__B2 _09688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10331_ _10331_/A _10331_/B vssd1 vssd1 vccd1 vccd1 _10331_/Y sky130_fd_sc_hd__nand2_1
XFILLER_139_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13050_ _18327_/Q _13046_/C _13049_/Y vssd1 vssd1 vccd1 vccd1 _18327_/D sky130_fd_sc_hd__o21a_1
X_10262_ _10262_/A _10262_/B vssd1 vssd1 vccd1 vccd1 _10262_/X sky130_fd_sc_hd__or2_1
XFILLER_152_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12001_ _17886_/A vssd1 vssd1 vccd1 vccd1 _12186_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17128__S _17130_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10193_ _09404_/A _10180_/X _10192_/X vssd1 vssd1 vccd1 vccd1 _10193_/X sky130_fd_sc_hd__a21o_1
XFILLER_78_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15300__A1 _15184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16967__S _16975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16740_ _16740_/A vssd1 vssd1 vccd1 vccd1 _16740_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13952_ _13769_/X _13773_/X _13968_/S vssd1 vssd1 vccd1 vccd1 _13952_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12903_ _18280_/Q _12910_/D _12933_/C vssd1 vssd1 vccd1 vccd1 _12907_/B sky130_fd_sc_hd__and3_1
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16671_ _19284_/Q _16670_/X _16671_/S vssd1 vssd1 vccd1 vccd1 _16672_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13883_ _13878_/X _13881_/X _14085_/S vssd1 vssd1 vccd1 vccd1 _13883_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18410_ _19788_/CLK _18410_/D vssd1 vssd1 vccd1 vccd1 _18410_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15172__A _15239_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15622_ _15622_/A vssd1 vssd1 vccd1 vccd1 _18829_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12834_ _12844_/A _12840_/C vssd1 vssd1 vccd1 vccd1 _12834_/Y sky130_fd_sc_hd__nor2_1
X_19390_ _19584_/CLK _19390_/D vssd1 vssd1 vccd1 vccd1 _19390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _19082_/CLK _18341_/D vssd1 vssd1 vccd1 vccd1 _18341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15553_/A vssd1 vssd1 vccd1 vccd1 _18804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _12765_/A _12810_/A vssd1 vssd1 vccd1 vccd1 _12765_/X sky130_fd_sc_hd__or2_1
XFILLER_15_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09294__A1 _18574_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14504_ _18225_/A vssd1 vssd1 vccd1 vccd1 _17862_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_125_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10523__S1 _10238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11205__A _11205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18272_ _19472_/CLK _18272_/D vssd1 vssd1 vccd1 vccd1 _18272_/Q sky130_fd_sc_hd__dfxtp_1
X_11716_ _11716_/A _11723_/B vssd1 vssd1 vccd1 vccd1 _11822_/D sky130_fd_sc_hd__nand2_2
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _15484_/A vssd1 vssd1 vccd1 vccd1 _18783_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12696_/A _16211_/B vssd1 vssd1 vccd1 vccd1 _12714_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17223_ _19493_/Q _17222_/X _17223_/S vssd1 vssd1 vccd1 vccd1 _17224_/A sky130_fd_sc_hd__mux2_1
X_14435_ _18490_/Q _19728_/Q _14443_/S vssd1 vssd1 vccd1 vccd1 _14436_/A sky130_fd_sc_hd__mux2_1
X_11647_ _12173_/A _11638_/Y _11646_/X vssd1 vssd1 vccd1 vccd1 _13650_/A sky130_fd_sc_hd__a21oi_4
XFILLER_168_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12478__A_N _12472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16207__S _16209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput13 io_dbus_rdata[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17154_ _10810_/X _13182_/X _17167_/S vssd1 vssd1 vccd1 vccd1 _17154_/X sky130_fd_sc_hd__mux2_1
Xinput24 io_dbus_rdata[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_2
XANTENNA__10287__S0 _09342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput35 io_ibus_inst[10] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15119__B2 _10098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14366_ _18467_/Q vssd1 vssd1 vccd1 vccd1 _14366_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput46 io_ibus_inst[20] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_2
X_11578_ _11501_/B _11528_/B _11339_/X vssd1 vssd1 vccd1 vccd1 _13573_/B sky130_fd_sc_hd__o21a_1
Xinput57 io_ibus_inst[30] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_2
XFILLER_155_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16105_ _16105_/A vssd1 vssd1 vccd1 vccd1 _19035_/D sky130_fd_sc_hd__clkbuf_1
Xinput68 io_irq_m2_irq vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__buf_8
X_13317_ _14514_/A vssd1 vssd1 vccd1 vccd1 _13317_/X sky130_fd_sc_hd__buf_2
XFILLER_155_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17085_ _17085_/A vssd1 vssd1 vccd1 vccd1 _19443_/D sky130_fd_sc_hd__clkbuf_1
X_10529_ _19511_/Q _19125_/Q _19575_/Q _18731_/Q _10558_/S _10367_/A vssd1 vssd1 vccd1
+ vccd1 _10530_/B sky130_fd_sc_hd__mux4_1
XFILLER_115_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14297_ _14297_/A _14300_/A vssd1 vssd1 vccd1 vccd1 _14297_/X sky130_fd_sc_hd__or2_1
XANTENNA__16731__A _16731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16036_ _16135_/S vssd1 vssd1 vccd1 vccd1 _16049_/S sky130_fd_sc_hd__buf_2
X_13248_ _13248_/A _18629_/Q vssd1 vssd1 vccd1 vccd1 _13248_/Y sky130_fd_sc_hd__nand2_1
XFILLER_112_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17816__A0 _15184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13179_ _12982_/B _13178_/X _12753_/A _19764_/Q vssd1 vssd1 vccd1 vccd1 _13179_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17987_ _19780_/Q _17988_/C _19781_/Q vssd1 vssd1 vccd1 vccd1 _17989_/B sky130_fd_sc_hd__a21oi_1
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19726_ _19726_/CLK _19726_/D vssd1 vssd1 vccd1 vccd1 _19726_/Q sky130_fd_sc_hd__dfxtp_1
X_16938_ _16768_/X _19378_/Q _16942_/S vssd1 vssd1 vccd1 vccd1 _16939_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10211__S0 _10094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19657_ _19657_/CLK _19657_/D vssd1 vssd1 vccd1 vccd1 _19657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16869_ _19348_/Q _16670_/X _16869_/S vssd1 vssd1 vccd1 vccd1 _16870_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10003__B _10003_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09410_ _10219_/A vssd1 vssd1 vccd1 vccd1 _09411_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18608_ _19329_/CLK _18608_/D vssd1 vssd1 vccd1 vccd1 _18608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19588_ _19589_/CLK _19588_/D vssd1 vssd1 vccd1 vccd1 _19588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10419__A1 _09171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09341_ _10277_/S vssd1 vssd1 vccd1 vccd1 _09342_/A sky130_fd_sc_hd__clkbuf_4
X_18539_ _18578_/CLK _18539_/D vssd1 vssd1 vccd1 vccd1 _18539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17501__S _17507_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15810__A _15878_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15358__A1 _15162_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09272_ _10857_/A _11046_/B vssd1 vssd1 vccd1 vccd1 _09273_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16117__S _16129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16641__A _16722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14333__A2 _12446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10658__A1 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09608_ _10325_/A vssd1 vssd1 vccd1 vccd1 _10177_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15597__A1 _15494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10880_ _18431_/Q _09280_/A _10857_/X _10879_/X vssd1 vssd1 vccd1 vccd1 _11779_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09539_ _09539_/A vssd1 vssd1 vccd1 vccd1 _09554_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11607__B1 _11602_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17411__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12550_ _12628_/A vssd1 vssd1 vccd1 vccd1 _12666_/B sky130_fd_sc_hd__buf_2
XANTENNA__15349__A1 _15149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11501_ _11551_/A _11501_/B vssd1 vssd1 vccd1 vccd1 _11664_/A sky130_fd_sc_hd__nand2_2
X_12481_ _12481_/A _12483_/B vssd1 vssd1 vccd1 vccd1 _12481_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16027__S _16027_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14220_ _14328_/A _14220_/B vssd1 vssd1 vccd1 vccd1 _14220_/Y sky130_fd_sc_hd__nand2_1
X_11432_ _11428_/Y _12765_/A _11430_/X _14582_/A vssd1 vssd1 vccd1 vccd1 _11432_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_172_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15866__S _15874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ _14155_/A _14155_/B vssd1 vssd1 vccd1 vccd1 _14151_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10075__S _10075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11363_ _11478_/A _11598_/B vssd1 vssd1 vccd1 vccd1 _11366_/B sky130_fd_sc_hd__nor2_1
XFILLER_153_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13102_ _17781_/A vssd1 vssd1 vccd1 vccd1 _13102_/X sky130_fd_sc_hd__buf_2
XFILLER_152_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10314_ _18601_/Q _19290_/Q _11156_/S vssd1 vssd1 vccd1 vccd1 _10314_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14082_ _14054_/X _14072_/X _14081_/Y _13784_/X vssd1 vssd1 vccd1 vccd1 _14082_/X
+ sky130_fd_sc_hd__o211a_1
X_11294_ _18557_/Q vssd1 vssd1 vccd1 vccd1 _14513_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_79_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17910_ _17910_/A vssd1 vssd1 vccd1 vccd1 _19757_/D sky130_fd_sc_hd__clkbuf_1
X_13033_ _13033_/A _18323_/Q _13033_/C vssd1 vssd1 vccd1 vccd1 _13034_/C sky130_fd_sc_hd__and3_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10245_ _10245_/A vssd1 vssd1 vccd1 vccd1 _10245_/X sky130_fd_sc_hd__buf_2
XFILLER_133_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18890_ _19444_/CLK _18890_/D vssd1 vssd1 vccd1 vccd1 _18890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10346__B1 _09625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17841_ _15219_/X _19721_/Q _17849_/S vssd1 vssd1 vccd1 vccd1 _17842_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10441__S0 _10230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ _19519_/Q _19133_/Q _19583_/Q _18739_/Q _09721_/X _09723_/X vssd1 vssd1 vccd1
+ vccd1 _10177_/B sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_51_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16697__S _16703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13296__C1 _13282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17772_ _19690_/Q _17771_/X _17772_/S vssd1 vssd1 vccd1 vccd1 _17773_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14984_ _14980_/X _14982_/Y _14983_/Y vssd1 vssd1 vccd1 vccd1 _16715_/A sky130_fd_sc_hd__a21oi_4
X_19511_ _19639_/CLK _19511_/D vssd1 vssd1 vccd1 vccd1 _19511_/Q sky130_fd_sc_hd__dfxtp_1
X_16723_ _19300_/Q _16721_/X _16735_/S vssd1 vssd1 vccd1 vccd1 _16724_/A sky130_fd_sc_hd__mux2_1
X_13935_ _10810_/X _13736_/X _13932_/X _13934_/Y vssd1 vssd1 vccd1 vccd1 _18430_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_81_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19442_ _19442_/CLK _19442_/D vssd1 vssd1 vccd1 vccd1 _19442_/Q sky130_fd_sc_hd__dfxtp_1
X_16654_ _16654_/A vssd1 vssd1 vccd1 vccd1 _16654_/X sky130_fd_sc_hd__clkbuf_2
X_13866_ _13745_/X _13665_/X _13806_/A vssd1 vssd1 vccd1 vccd1 _13866_/X sky130_fd_sc_hd__a21o_1
X_15605_ _15662_/S vssd1 vssd1 vccd1 vccd1 _15614_/S sky130_fd_sc_hd__buf_2
XFILLER_34_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12817_ _18173_/A vssd1 vssd1 vccd1 vccd1 _12817_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13134__B _13134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19373_ _19537_/CLK _19373_/D vssd1 vssd1 vccd1 vccd1 _19373_/Q sky130_fd_sc_hd__dfxtp_1
X_16585_ _19248_/Q vssd1 vssd1 vccd1 vccd1 _16586_/A sky130_fd_sc_hd__clkbuf_1
X_13797_ _13797_/A vssd1 vssd1 vccd1 vccd1 _13797_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18324_ _18330_/CLK _18324_/D vssd1 vssd1 vccd1 vccd1 _18324_/Q sky130_fd_sc_hd__dfxtp_1
X_15536_ _18799_/Q _15535_/X _15536_/S vssd1 vssd1 vccd1 vccd1 _15537_/A sky130_fd_sc_hd__mux2_1
X_12748_ _12748_/A vssd1 vssd1 vccd1 vccd1 _12749_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11074__B2 _12466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18255_ _19855_/CLK _18255_/D vssd1 vssd1 vccd1 vccd1 _18255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15467_ _15467_/A vssd1 vssd1 vccd1 vccd1 _18775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12679_ _19662_/Q _12668_/X _12672_/X _12678_/X vssd1 vssd1 vccd1 vccd1 _12679_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17206_ _19488_/Q _17205_/X _17206_/S vssd1 vssd1 vccd1 vccd1 _17207_/A sky130_fd_sc_hd__mux2_1
X_14418_ _18485_/Q vssd1 vssd1 vccd1 vccd1 _15027_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18186_ _18197_/A _18191_/C vssd1 vssd1 vccd1 vccd1 _18186_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15398_ _18746_/Q _15219_/X _15406_/S vssd1 vssd1 vccd1 vccd1 _15399_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17137_ _11463_/B _11463_/C _11822_/D vssd1 vssd1 vccd1 vccd1 _17137_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15776__S _15780_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14349_ _17621_/A _18493_/Q _14352_/S vssd1 vssd1 vccd1 vccd1 _14350_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_1_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_6_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17068_ _17068_/A vssd1 vssd1 vccd1 vccd1 _19435_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16019_ _15009_/X _19007_/Q _16027_/S vssd1 vssd1 vccd1 vccd1 _16020_/A sky130_fd_sc_hd__mux2_1
X_09890_ _09942_/A _09890_/B vssd1 vssd1 vccd1 vccd1 _09890_/Y sky130_fd_sc_hd__nor2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10888__A1 _09353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16400__S _16402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09803__A _09803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19709_ _19709_/CLK _19709_/D vssd1 vssd1 vccd1 vccd1 _19709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11544__S _14032_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14251__A1 _14126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ _10850_/A vssd1 vssd1 vccd1 vccd1 _10640_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_167_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10499__S0 _10242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12793__A_N _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11160__S1 _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10273__C1 _09248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09255_ _09255_/A vssd1 vssd1 vccd1 vccd1 _16212_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_166_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17740__A2 _12779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09186_ _10210_/A vssd1 vssd1 vccd1 vccd1 _10107_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_135_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_162_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19692_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_88_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16371__A _16428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12317__A1 _19684_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09718__C1 _09708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_177_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19703_/CLK sky130_fd_sc_hd__clkbuf_16
X_10030_ _19264_/Q _19035_/Q _18966_/Q _19360_/Q _09952_/S _10029_/X vssd1 vssd1 vccd1
+ vccd1 _10030_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10423__S0 _11088_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10879__B2 _10823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10974__S1 _10906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16310__S _16318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_3_0_clock clkbuf_4_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_100_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _18395_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11981_ _19736_/Q _19737_/Q _19738_/Q _19739_/Q vssd1 vssd1 vccd1 vccd1 _12093_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__14490__A1 _19753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13235__A _13235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13720_ _13720_/A _13720_/B _13922_/A vssd1 vssd1 vccd1 vccd1 _14003_/A sky130_fd_sc_hd__nor3_2
X_10932_ _18852_/Q _19310_/Q _10932_/S vssd1 vssd1 vccd1 vccd1 _10933_/B sky130_fd_sc_hd__mux2_1
XFILLER_72_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13651_ _13993_/A vssd1 vssd1 vccd1 vccd1 _13968_/S sky130_fd_sc_hd__clkbuf_2
X_10863_ _10873_/A _10863_/B vssd1 vssd1 vccd1 vccd1 _10863_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_115_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _18564_/CLK sky130_fd_sc_hd__clkbuf_16
X_12602_ _12602_/A vssd1 vssd1 vccd1 vccd1 _12602_/X sky130_fd_sc_hd__buf_2
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _16370_/A vssd1 vssd1 vccd1 vccd1 _19151_/D sky130_fd_sc_hd__clkbuf_1
X_13582_ _13720_/A _13785_/A vssd1 vssd1 vccd1 vccd1 _13783_/B sky130_fd_sc_hd__nor2_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ _18757_/Q _18986_/Q _18917_/Q _19215_/Q _10934_/S _10785_/A vssd1 vssd1 vccd1
+ vccd1 _10795_/B sky130_fd_sc_hd__mux4_1
XFILLER_9_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _15321_/A vssd1 vssd1 vccd1 vccd1 _18712_/D sky130_fd_sc_hd__clkbuf_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10264__C1 _09134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12533_ _12533_/A _12533_/B _12540_/A vssd1 vssd1 vccd1 vccd1 _12751_/C sky130_fd_sc_hd__or3_2
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16980__S _16986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17731__A2 _13346_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18040_ _18043_/A _18043_/C _18039_/X vssd1 vssd1 vccd1 vccd1 _18040_/Y sky130_fd_sc_hd__a21oi_1
X_15252_ _18685_/Q _15251_/X _15260_/S vssd1 vssd1 vccd1 vccd1 _15253_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12464_ _12464_/A vssd1 vssd1 vccd1 vccd1 _12464_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14203_ _14203_/A _14203_/B vssd1 vssd1 vccd1 vccd1 _14203_/Y sky130_fd_sc_hd__nor2_1
X_11415_ _18542_/Q vssd1 vssd1 vccd1 vccd1 _11821_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11202__B _12504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15183_ _15183_/A vssd1 vssd1 vccd1 vccd1 _18664_/D sky130_fd_sc_hd__clkbuf_1
X_12395_ _19756_/Q _12116_/X _12391_/X _12394_/Y vssd1 vssd1 vccd1 vccd1 _17907_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_125_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09594__S _10185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14134_ _18440_/Q _14120_/X _14133_/X vssd1 vssd1 vccd1 vccd1 _18440_/D sky130_fd_sc_hd__o21a_1
XFILLER_153_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11346_ _11346_/A vssd1 vssd1 vccd1 vccd1 _11642_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14513__B _14519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09709__C1 _09708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14065_ _14314_/A _14220_/B vssd1 vssd1 vccd1 vccd1 _14065_/Y sky130_fd_sc_hd__nor2_1
X_18942_ _19592_/CLK _18942_/D vssd1 vssd1 vccd1 vccd1 _18942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12314__A _19753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ _11225_/X _11226_/Y _11274_/X _11275_/Y _11276_/Y vssd1 vssd1 vccd1 vccd1
+ _11277_/X sky130_fd_sc_hd__o2111a_1
X_13016_ _13034_/A _13016_/B _13016_/C vssd1 vssd1 vccd1 vccd1 _18317_/D sky130_fd_sc_hd__nor3_1
X_10228_ _19518_/Q _19132_/Q _19582_/Q _18738_/Q _09583_/A _10390_/A vssd1 vssd1 vccd1
+ vccd1 _10229_/B sky130_fd_sc_hd__mux4_2
X_18873_ _19331_/CLK _18873_/D vssd1 vssd1 vccd1 vccd1 _18873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17824_ _17824_/A vssd1 vssd1 vccd1 vccd1 _19713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__16220__S _16224_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10159_ _10212_/A _10159_/B vssd1 vssd1 vccd1 vccd1 _10159_/X sky130_fd_sc_hd__or2_1
XFILLER_67_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17755_ _19686_/Q _17708_/A _17753_/Y _17754_/X vssd1 vssd1 vccd1 vccd1 _19686_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14967_ _17728_/A _14979_/C vssd1 vssd1 vccd1 vccd1 _14969_/B sky130_fd_sc_hd__nor2_1
XANTENNA__14481__A1 _19749_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16706_ _16722_/A vssd1 vssd1 vccd1 vccd1 _16719_/S sky130_fd_sc_hd__buf_4
XANTENNA__17840__A _17840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13918_ _13915_/X _13917_/X _13918_/S vssd1 vssd1 vccd1 vccd1 _13918_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17686_ _13307_/X _17685_/Y _17686_/S vssd1 vssd1 vccd1 vccd1 _17686_/X sky130_fd_sc_hd__mux2_1
X_14898_ _19080_/Q vssd1 vssd1 vccd1 vccd1 _14898_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19425_ _19838_/CLK _19425_/D vssd1 vssd1 vccd1 vccd1 _19425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16637_ _19274_/Q vssd1 vssd1 vccd1 vccd1 _16638_/A sky130_fd_sc_hd__clkbuf_1
X_13849_ _13812_/X _13848_/Y _13997_/S vssd1 vssd1 vccd1 vccd1 _13946_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19356_ _19613_/CLK _19356_/D vssd1 vssd1 vccd1 vccd1 _19356_/Q sky130_fd_sc_hd__dfxtp_1
X_16568_ _16568_/A vssd1 vssd1 vccd1 vccd1 _19239_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18307_ _18329_/CLK _18307_/D vssd1 vssd1 vccd1 vccd1 _18307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15519_ _16774_/A vssd1 vssd1 vccd1 vccd1 _15519_/X sky130_fd_sc_hd__clkbuf_2
X_16499_ _16131_/X _19209_/Q _16501_/S vssd1 vssd1 vccd1 vccd1 _16500_/A sky130_fd_sc_hd__mux2_1
X_19287_ _19546_/CLK _19287_/D vssd1 vssd1 vccd1 vccd1 _19287_/Q sky130_fd_sc_hd__dfxtp_1
X_18238_ _18239_/B _18239_/C _18237_/Y vssd1 vssd1 vccd1 vccd1 _19867_/D sky130_fd_sc_hd__o21a_1
XANTENNA__12208__B _14216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18169_ _19843_/Q _18167_/B _18168_/Y vssd1 vssd1 vccd1 vccd1 _19843_/D sky130_fd_sc_hd__o21a_1
XFILLER_144_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10653__S0 _10500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13523__D_N _11517_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_94_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19858_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09942_ _09942_/A _09942_/B vssd1 vssd1 vccd1 vccd1 _09942_/X sky130_fd_sc_hd__or2_1
XFILLER_143_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17238__A1 _13412_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09873_ _09873_/A vssd1 vssd1 vccd1 vccd1 _09873_/Y sky130_fd_sc_hd__inv_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15535__A _16790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11782__B _13630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15254__B _15254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14472__A1 _19745_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_32_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19553_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12894__A _12904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09307_ _09307_/A vssd1 vssd1 vccd1 vccd1 _09308_/A sky130_fd_sc_hd__buf_2
XFILLER_166_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19331_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17174__A0 _18436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09238_ _18848_/Q _19402_/Q _19564_/Q _18816_/Q _09190_/X _09165_/A vssd1 vssd1 vccd1
+ vccd1 _09238_/X sky130_fd_sc_hd__mux4_1
XANTENNA__14527__A2 _12763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17909__B _17909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09169_ _09169_/A vssd1 vssd1 vccd1 vccd1 _09170_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ _11200_/A _12503_/A vssd1 vssd1 vccd1 vccd1 _11251_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09708__A _09708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10644__S0 _10631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12180_ _12180_/A vssd1 vssd1 vccd1 vccd1 _14203_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11761__A2 _11022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ _11131_/A _11130_/Y vssd1 vssd1 vccd1 vccd1 _11132_/A sky130_fd_sc_hd__or2b_1
XANTENNA__17925__A _19760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17229__A1 _13376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11062_ _11062_/A _11062_/B vssd1 vssd1 vccd1 vccd1 _11062_/X sky130_fd_sc_hd__or2_1
XFILLER_77_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17136__S _17143_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ _09783_/X _10010_/X _10012_/X vssd1 vssd1 vccd1 vccd1 _10013_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10947__S1 _10772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15870_ _15033_/X _18940_/Q _15874_/S vssd1 vssd1 vccd1 vccd1 _15871_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16040__S _16049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A io_dbus_rdata[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ _16774_/A vssd1 vssd1 vccd1 vccd1 _14821_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16975__S _16975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10589__A _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14463__A1 _12043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14752_ _16651_/A vssd1 vssd1 vccd1 vccd1 _16755_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17540_ _19630_/Q _16749_/A _17546_/S vssd1 vssd1 vccd1 vccd1 _17541_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11964_ _11885_/X _11961_/X _11963_/Y _11625_/A vssd1 vssd1 vccd1 vccd1 _11964_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09565__S1 _09144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13703_ _13703_/A vssd1 vssd1 vccd1 vccd1 _13818_/B sky130_fd_sc_hd__clkbuf_2
X_17471_ _17471_/A vssd1 vssd1 vccd1 vccd1 _19599_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10915_ _19693_/Q _10915_/B vssd1 vssd1 vccd1 vccd1 _10915_/X sky130_fd_sc_hd__or2_1
X_14683_ _14683_/A vssd1 vssd1 vccd1 vccd1 _18580_/D sky130_fd_sc_hd__clkbuf_1
X_11895_ _14045_/A _11895_/B vssd1 vssd1 vccd1 vccd1 _11922_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__10101__B _12489_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output109_A _12495_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11029__A1 _09169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19210_ _19727_/CLK _19210_/D vssd1 vssd1 vccd1 vccd1 _19210_/Q sky130_fd_sc_hd__dfxtp_1
X_16422_ _19175_/Q _15580_/X _16424_/S vssd1 vssd1 vccd1 vccd1 _16423_/A sky130_fd_sc_hd__mux2_1
X_13634_ _13765_/S vssd1 vssd1 vccd1 vccd1 _13741_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_44_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10846_ _10846_/A _10846_/B _10846_/C vssd1 vssd1 vccd1 vccd1 _10846_/X sky130_fd_sc_hd__or3_2
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11124__S1 _10245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19141_ _19622_/CLK _19141_/D vssd1 vssd1 vccd1 vccd1 _19141_/Q sky130_fd_sc_hd__dfxtp_1
X_16353_ _16131_/X _19145_/Q _16355_/S vssd1 vssd1 vccd1 vccd1 _16354_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13565_ _15095_/A vssd1 vssd1 vccd1 vccd1 _15116_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_158_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10777_ _18759_/Q _18988_/Q _18919_/Q _19217_/Q _10934_/S _10713_/A vssd1 vssd1 vccd1
+ vccd1 _10778_/B sky130_fd_sc_hd__mux4_2
X_15304_ _15304_/A vssd1 vssd1 vccd1 vccd1 _18704_/D sky130_fd_sc_hd__clkbuf_1
X_12516_ _12516_/A vssd1 vssd1 vccd1 vccd1 _12664_/A sky130_fd_sc_hd__clkbuf_2
X_19072_ _19622_/CLK _19072_/D vssd1 vssd1 vccd1 vccd1 _19072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16284_ _16284_/A vssd1 vssd1 vccd1 vccd1 _19114_/D sky130_fd_sc_hd__clkbuf_1
X_13496_ _13496_/A vssd1 vssd1 vccd1 vccd1 _18406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18023_ _18023_/A _18023_/B _19794_/Q vssd1 vssd1 vccd1 vccd1 _18025_/B sky130_fd_sc_hd__and3_1
X_15235_ _16737_/A vssd1 vssd1 vccd1 vccd1 _15235_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12447_ _14331_/A _12447_/B vssd1 vssd1 vccd1 vccd1 _13590_/S sky130_fd_sc_hd__nand2_2
XFILLER_138_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output90_A _12313_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10635__S0 _10631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15166_ _18659_/Q _15165_/X _15169_/S vssd1 vssd1 vccd1 vccd1 _15167_/A sky130_fd_sc_hd__mux2_1
X_12378_ _13712_/A _14289_/A _12350_/B vssd1 vssd1 vccd1 vccd1 _12379_/B sky130_fd_sc_hd__a21oi_1
XFILLER_114_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14117_ _12013_/X _14102_/X _14116_/X vssd1 vssd1 vccd1 vccd1 _14117_/X sky130_fd_sc_hd__a21bo_1
XFILLER_113_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11329_ _11375_/B _11640_/B vssd1 vssd1 vccd1 vccd1 _11584_/B sky130_fd_sc_hd__nor2_1
XFILLER_125_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12044__A _12067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15097_ _15111_/A vssd1 vssd1 vccd1 vccd1 _15097_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_141_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18925_ _19223_/CLK _18925_/D vssd1 vssd1 vccd1 vccd1 _18925_/Q sky130_fd_sc_hd__dfxtp_1
X_14048_ _14037_/X _14038_/Y _14047_/X _13594_/A vssd1 vssd1 vccd1 vccd1 _14048_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10938__S1 _09352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18856_ _19569_/CLK _18856_/D vssd1 vssd1 vccd1 vccd1 _18856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09353__A _09353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17807_ _17853_/S vssd1 vssd1 vccd1 vccd1 _17816_/S sky130_fd_sc_hd__buf_4
XFILLER_83_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18787_ _19537_/CLK _18787_/D vssd1 vssd1 vccd1 vccd1 _18787_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14454__A1 _19737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16885__S _16891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15999_ _14908_/X _18998_/Q _16005_/S vssd1 vssd1 vccd1 vccd1 _16000_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17570__A _17592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17738_ _17737_/A _17737_/C _14990_/A vssd1 vssd1 vccd1 vccd1 _17738_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09556__S1 _09555_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17669_ _17674_/B _17669_/B vssd1 vssd1 vccd1 vccd1 _17669_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13603__A _13603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19408_ _19506_/CLK _19408_/D vssd1 vssd1 vccd1 vccd1 _19408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13414__C1 _13401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19339_ _19632_/CLK _19339_/D vssd1 vssd1 vccd1 vccd1 _19339_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_173_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11123__A _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10874__S0 _10614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15964__S _15972_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09925_ _09925_/A vssd1 vssd1 vccd1 vccd1 _09926_/A sky130_fd_sc_hd__buf_2
XFILLER_59_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14595__A2_N _12731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14693__A1 _14587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13484__S _13486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14693__B2 input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09856_ _09856_/A _09856_/B vssd1 vssd1 vccd1 vccd1 _09856_/X sky130_fd_sc_hd__or2_1
XFILLER_131_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10703__B1 _10793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_98_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09787_ _19653_/Q _19070_/Q _19107_/Q _18713_/Q _09760_/X _09763_/X vssd1 vssd1 vccd1
+ vccd1 _09788_/B sky130_fd_sc_hd__mux4_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16795__S _16807_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _19604_/Q _19442_/Q _18888_/Q _18658_/Q _10886_/S _09352_/A vssd1 vssd1 vccd1
+ vccd1 _10701_/B sky130_fd_sc_hd__mux4_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13405__C1 _13404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11680_ _16212_/D vssd1 vssd1 vccd1 vccd1 _11994_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11106__S1 _10245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ _10631_/A vssd1 vssd1 vccd1 vccd1 _10631_/X sky130_fd_sc_hd__buf_4
XFILLER_139_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10348__S _10348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13350_ _14514_/A vssd1 vssd1 vccd1 vccd1 _13350_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10865__S0 _09152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10562_ _19252_/Q _19023_/Q _18954_/Q _19348_/Q _10540_/S _09141_/A vssd1 vssd1 vccd1
+ vccd1 _10562_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12301_ _12296_/Y _12300_/X _19752_/Q _12002_/X vssd1 vssd1 vccd1 vccd1 _12301_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_127_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13281_ _17892_/A vssd1 vssd1 vccd1 vccd1 _14514_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10493_ _10498_/A _10490_/X _10492_/X _09681_/A vssd1 vssd1 vccd1 vccd1 _10494_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13184__A1 _13139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15020_ _14711_/X _15013_/Y _15019_/X vssd1 vssd1 vccd1 vccd1 _16725_/A sky130_fd_sc_hd__o21ai_4
X_12232_ _10003_/B _12328_/A _12231_/X vssd1 vssd1 vccd1 vccd1 _13615_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__10617__S0 _10614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15874__S _15874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12163_ _12163_/A _12163_/B vssd1 vssd1 vccd1 vccd1 _12163_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__09872__S _09872_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11114_ _19256_/Q _19027_/Q _18958_/Q _19352_/Q _11110_/S _09483_/X vssd1 vssd1 vccd1
+ vccd1 _11114_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16971_ _16816_/X _19393_/Q _16975_/S vssd1 vssd1 vccd1 vccd1 _16972_/A sky130_fd_sc_hd__mux2_1
X_12094_ _19734_/Q _19735_/Q _19743_/Q _12094_/D vssd1 vssd1 vccd1 vccd1 _12117_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14684__A1 _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18710_ _19618_/CLK _18710_/D vssd1 vssd1 vccd1 vccd1 _18710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14684__B2 input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15175__A _16677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11042__S0 _10919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11045_ _18426_/Q vssd1 vssd1 vccd1 vccd1 _11046_/A sky130_fd_sc_hd__clkbuf_8
X_15922_ _14929_/X _18963_/Q _15924_/S vssd1 vssd1 vccd1 vccd1 _15923_/A sky130_fd_sc_hd__mux2_1
X_19690_ _19690_/CLK _19690_/D vssd1 vssd1 vccd1 vccd1 _19690_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_103_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09173__A _09173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18641_ _19628_/CLK _18641_/D vssd1 vssd1 vccd1 vccd1 _18641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15853_ _15853_/A vssd1 vssd1 vccd1 vccd1 _18932_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13239__A2 _12668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_0_0_clock clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_64_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14804_ _14804_/A vssd1 vssd1 vccd1 vccd1 _14804_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18572_ _18578_/CLK _18572_/D vssd1 vssd1 vccd1 vccd1 _18572_/Q sky130_fd_sc_hd__dfxtp_1
X_12996_ _13006_/D vssd1 vssd1 vccd1 vccd1 _13003_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15784_ _15784_/A vssd1 vssd1 vccd1 vccd1 _18901_/D sky130_fd_sc_hd__clkbuf_1
X_17523_ _19623_/Q _16725_/X _17529_/S vssd1 vssd1 vccd1 vccd1 _17524_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11947_ _11947_/A _14075_/B vssd1 vssd1 vccd1 vccd1 _11953_/A sky130_fd_sc_hd__xor2_1
X_14735_ _18428_/Q _14958_/A _14875_/A vssd1 vssd1 vccd1 vccd1 _14735_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09863__A1 _09217_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ _17454_/A vssd1 vssd1 vccd1 vccd1 _19592_/D sky130_fd_sc_hd__clkbuf_1
X_14666_ _14677_/A _15954_/B vssd1 vssd1 vccd1 vccd1 _14667_/A sky130_fd_sc_hd__and2_1
X_11878_ _11844_/B _11873_/X _11877_/X vssd1 vssd1 vccd1 vccd1 _11879_/B sky130_fd_sc_hd__a21o_2
X_16405_ _19167_/Q _15554_/X _16413_/S vssd1 vssd1 vccd1 vccd1 _16406_/A sky130_fd_sc_hd__mux2_1
X_13617_ _13617_/A vssd1 vssd1 vccd1 vccd1 _14026_/B sky130_fd_sc_hd__clkbuf_2
X_10829_ _18821_/Q _19375_/Q _19537_/Q _18789_/Q _11027_/S _10813_/A vssd1 vssd1 vccd1
+ vccd1 _10830_/B sky130_fd_sc_hd__mux4_1
XANTENNA__14953__S _14997_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14597_ _18205_/A vssd1 vssd1 vccd1 vccd1 _14597_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17385_ _16838_/X _19562_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _17386_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16734__A _16734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19124_ _19713_/CLK _19124_/D vssd1 vssd1 vccd1 vccd1 _19124_/Q sky130_fd_sc_hd__dfxtp_1
X_16336_ _16106_/X _19137_/Q _16340_/S vssd1 vssd1 vccd1 vccd1 _16337_/A sky130_fd_sc_hd__mux2_1
X_13548_ _13560_/A _13548_/B vssd1 vssd1 vccd1 vccd1 _13549_/A sky130_fd_sc_hd__and2_1
XFILLER_118_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16267_ _16267_/A vssd1 vssd1 vccd1 vccd1 _19106_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19055_ _19712_/CLK _19055_/D vssd1 vssd1 vccd1 vccd1 _19055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13479_ _13479_/A vssd1 vssd1 vccd1 vccd1 _18398_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16361__A1 _15487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15218_ _15218_/A vssd1 vssd1 vccd1 vccd1 _18675_/D sky130_fd_sc_hd__clkbuf_1
X_18006_ hold2/X _19786_/Q _18006_/C vssd1 vssd1 vccd1 vccd1 _18011_/C sky130_fd_sc_hd__and3_1
XANTENNA__09348__A _09928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16198_ _16198_/A vssd1 vssd1 vccd1 vccd1 _19071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10528__A3 _10527_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15149_ _16651_/A vssd1 vssd1 vccd1 vccd1 _15149_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_141_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09710_ _09689_/X _09694_/X _09703_/X _09709_/X _09134_/A vssd1 vssd1 vccd1 vccd1
+ _09710_/X sky130_fd_sc_hd__a311o_2
XFILLER_68_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18908_ _19592_/CLK _18908_/D vssd1 vssd1 vccd1 vccd1 _18908_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09777__S1 _09763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__A _12502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09641_ _18613_/Q _19302_/Q _10417_/S vssd1 vssd1 vccd1 vccd1 _09642_/B sky130_fd_sc_hd__mux2_1
X_18839_ _19587_/CLK _18839_/D vssd1 vssd1 vccd1 vccd1 _18839_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10161__A1 _10007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09572_ _09772_/A _09569_/X _09571_/X _09562_/X vssd1 vssd1 vccd1 vccd1 _09572_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09606__A1 _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13402__A2 _13399_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10847__S0 _10648_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11788__A _19733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14164__A _14168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12913__A1 _18282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09908_ _09908_/A _09908_/B vssd1 vssd1 vccd1 vccd1 _09908_/X sky130_fd_sc_hd__or2_1
XANTENNA__12412__A _19688_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09839_ _09430_/X _09817_/X _09837_/X _09625_/X _09838_/Y vssd1 vssd1 vccd1 vccd1
+ _12497_/A sky130_fd_sc_hd__o32a_4
XFILLER_46_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16819__A _16819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12850_ _18265_/Q _12850_/B _12850_/C vssd1 vssd1 vccd1 vccd1 _12851_/C sky130_fd_sc_hd__and3_1
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _11801_/A vssd1 vssd1 vccd1 vccd1 _11801_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _18302_/Q _12780_/X _16211_/B vssd1 vssd1 vccd1 vccd1 _12781_/X sky130_fd_sc_hd__mux2_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09845__A1 _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _18527_/Q _12692_/X _14519_/X _14514_/X vssd1 vssd1 vccd1 vccd1 _18527_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11732_ _13653_/A _13996_/A vssd1 vssd1 vccd1 vccd1 _11733_/B sky130_fd_sc_hd__and2b_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14451_ _14451_/A vssd1 vssd1 vccd1 vccd1 _18497_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _11752_/C vssd1 vssd1 vccd1 vccd1 _11663_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13402_ _13354_/X _13399_/X _13400_/X _13401_/X vssd1 vssd1 vccd1 vccd1 _18378_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17170_ _17204_/A vssd1 vssd1 vccd1 vccd1 _17184_/S sky130_fd_sc_hd__clkbuf_2
X_10614_ _11028_/S vssd1 vssd1 vccd1 vccd1 _10614_/X sky130_fd_sc_hd__buf_4
X_14382_ _14382_/A vssd1 vssd1 vccd1 vccd1 _18472_/D sky130_fd_sc_hd__clkbuf_1
X_11594_ _12259_/B _12259_/C vssd1 vssd1 vccd1 vccd1 _11697_/S sky130_fd_sc_hd__nor2_4
X_16121_ _16121_/A vssd1 vssd1 vccd1 vccd1 _19040_/D sky130_fd_sc_hd__clkbuf_1
X_13333_ _18640_/Q _14958_/B _14958_/C _14958_/D vssd1 vssd1 vccd1 vccd1 _13333_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__10758__A3 _10757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10545_ _10910_/A vssd1 vssd1 vccd1 vccd1 _10739_/A sky130_fd_sc_hd__buf_2
XFILLER_155_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16052_ _16135_/S vssd1 vssd1 vccd1 vccd1 _16065_/S sky130_fd_sc_hd__buf_2
X_13264_ _12713_/X _13118_/X _13263_/X _13232_/X vssd1 vssd1 vccd1 vccd1 _18361_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10476_ _19512_/Q _19126_/Q _19576_/Q _18732_/Q _09631_/A _10368_/A vssd1 vssd1 vccd1
+ vccd1 _10477_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12365__C1 _12193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15003_ _14990_/A _15002_/C _18483_/Q vssd1 vssd1 vccd1 vccd1 _15003_/Y sky130_fd_sc_hd__a21oi_1
X_12215_ _19747_/Q _19748_/Q _12215_/C vssd1 vssd1 vccd1 vccd1 _12217_/B sky130_fd_sc_hd__and3_1
XFILLER_29_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13195_ _17944_/B _13123_/A _13191_/X _13194_/X vssd1 vssd1 vccd1 vccd1 _13196_/B
+ sky130_fd_sc_hd__a211o_2
XANTENNA__10107__A _10107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19811_ _19812_/CLK _19811_/D vssd1 vssd1 vccd1 vccd1 _19811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12146_ _12142_/A _12145_/X _12411_/B vssd1 vssd1 vccd1 vccd1 _12146_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_121_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14657__A1 _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10391__A1 _10239_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14657__B2 input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19742_ _19753_/CLK _19742_/D vssd1 vssd1 vccd1 vccd1 _19742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12077_ _19743_/Q _11788_/B _12073_/X _12076_/Y vssd1 vssd1 vccd1 vccd1 _17884_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_110_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16954_ _16954_/A vssd1 vssd1 vccd1 vccd1 _19385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09533__B1 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15905_ _14833_/X _18955_/Q _15913_/S vssd1 vssd1 vccd1 vccd1 _15906_/A sky130_fd_sc_hd__mux2_1
X_11028_ _18849_/Q _19307_/Q _11028_/S vssd1 vssd1 vccd1 vccd1 _11028_/X sky130_fd_sc_hd__mux2_1
X_19673_ _19686_/CLK _19673_/D vssd1 vssd1 vccd1 vccd1 _19673_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16885_ _19355_/Q _16693_/X _16891_/S vssd1 vssd1 vccd1 vccd1 _16886_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18624_ _19692_/CLK _18624_/D vssd1 vssd1 vccd1 vccd1 _18624_/Q sky130_fd_sc_hd__dfxtp_2
X_15836_ _15836_/A vssd1 vssd1 vccd1 vccd1 _18924_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11891__B2 _11788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09631__A _09631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18555_ _18564_/CLK _18555_/D vssd1 vssd1 vccd1 vccd1 _18555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09836__A1 _09819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12979_ _12982_/B _12982_/C _12922_/X vssd1 vssd1 vccd1 vccd1 _12979_/Y sky130_fd_sc_hd__a21oi_1
X_15767_ _14867_/X _18894_/Q _15769_/S vssd1 vssd1 vccd1 vccd1 _15768_/A sky130_fd_sc_hd__mux2_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17506_ _17506_/A vssd1 vssd1 vccd1 vccd1 _19615_/D sky130_fd_sc_hd__clkbuf_1
X_14718_ _16212_/C _14718_/B vssd1 vssd1 vccd1 vccd1 _15960_/C sky130_fd_sc_hd__nand2_1
X_18486_ _19686_/CLK _18486_/D vssd1 vssd1 vccd1 vccd1 _18486_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15698_ _15698_/A vssd1 vssd1 vccd1 vccd1 _18863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17437_ _17448_/A vssd1 vssd1 vccd1 vccd1 _17446_/S sky130_fd_sc_hd__buf_4
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14649_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14649_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_46_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10829__S0 _11027_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17368_ _16813_/X _19554_/Q _17374_/S vssd1 vssd1 vccd1 vccd1 _17369_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19107_ _19718_/CLK _19107_/D vssd1 vssd1 vccd1 vccd1 _19107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16319_ _16319_/A vssd1 vssd1 vccd1 vccd1 _19129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17299_ _17299_/A vssd1 vssd1 vccd1 vccd1 _19523_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19038_ _19589_/CLK _19038_/D vssd1 vssd1 vccd1 vccd1 _19038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput101 _11813_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[6] sky130_fd_sc_hd__buf_2
Xoutput112 _12477_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[10] sky130_fd_sc_hd__buf_2
Xoutput123 _12490_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[20] sky130_fd_sc_hd__buf_2
XFILLER_126_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15808__A _17391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput134 _12504_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[30] sky130_fd_sc_hd__buf_2
Xoutput145 _17874_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[10] sky130_fd_sc_hd__buf_2
Xoutput156 _12201_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[20] sky130_fd_sc_hd__buf_2
XFILLER_115_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput167 _12441_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[30] sky130_fd_sc_hd__buf_2
XANTENNA__09806__A _09819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11174__A3 _11173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14431__B _14431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11006__S0 _10724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13320__A1 _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09624_ _09624_/A _09624_/B vssd1 vssd1 vccd1 vccd1 _09625_/A sky130_fd_sc_hd__nand2_4
XFILLER_55_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15073__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09541__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15262__B _15262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09555_ _09642_/A vssd1 vssd1 vccd1 vccd1 _09555_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11095__C1 _10373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09260__B _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09486_ _10384_/A vssd1 vssd1 vccd1 vccd1 _09486_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09460__C1 _09459_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12407__A _12408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10070__B1 _09318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10330_ _18601_/Q _19290_/Q _11188_/S vssd1 vssd1 vccd1 vccd1 _10331_/B sky130_fd_sc_hd__mux2_1
XFILLER_137_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17409__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ _18769_/Q _18998_/Q _18929_/Q _19227_/Q _09793_/A _09144_/A vssd1 vssd1 vccd1
+ vccd1 _10262_/B sky130_fd_sc_hd__mux4_1
XFILLER_106_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12000_ _12116_/A vssd1 vssd1 vccd1 vccd1 _17886_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10192_ _09621_/X _10182_/Y _10187_/X _10191_/Y _09395_/A vssd1 vssd1 vccd1 vccd1
+ _10192_/X sky130_fd_sc_hd__o311a_1
XFILLER_79_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12142__A _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13951_ _14130_/A _13944_/X _13949_/Y _13950_/X vssd1 vssd1 vccd1 vccd1 _13951_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13672__S _13724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ _12910_/D _12933_/C _18280_/Q vssd1 vssd1 vccd1 vccd1 _12904_/B sky130_fd_sc_hd__a21oi_1
X_13882_ _13969_/S vssd1 vssd1 vccd1 vccd1 _14085_/S sky130_fd_sc_hd__clkbuf_2
X_16670_ _16670_/A vssd1 vssd1 vccd1 vccd1 _16670_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15064__A1 _11542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12833_ _12842_/D vssd1 vssd1 vccd1 vccd1 _12840_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15621_ _18829_/Q _15529_/X _15625_/S vssd1 vssd1 vccd1 vccd1 _15622_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _18401_/CLK _18340_/D vssd1 vssd1 vccd1 vccd1 _18340_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _12731_/X _12732_/X _12759_/X _12763_/X vssd1 vssd1 vccd1 vccd1 _18299_/D
+ sky130_fd_sc_hd__o22a_1
X_15552_ _18804_/Q _15551_/X _15552_/S vssd1 vssd1 vccd1 vccd1 _15553_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _11821_/A _18299_/Q vssd1 vssd1 vccd1 vccd1 _11715_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10833__C1 _09244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15599__S _15603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14503_ _14503_/A vssd1 vssd1 vccd1 vccd1 _18521_/D sky130_fd_sc_hd__clkbuf_1
X_18271_ _19472_/CLK _18271_/D vssd1 vssd1 vccd1 vccd1 _18271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15483_ _18783_/Q _15235_/X _15485_/S vssd1 vssd1 vccd1 vccd1 _15484_/A sky130_fd_sc_hd__mux2_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11205__B _12505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12695_ _17882_/A vssd1 vssd1 vccd1 vccd1 _17774_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17222_ _18450_/Q _12779_/X _17235_/S vssd1 vssd1 vccd1 vccd1 _17222_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13701__A _13761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11646_ _12005_/A _12462_/A vssd1 vssd1 vccd1 vccd1 _11646_/X sky130_fd_sc_hd__and2b_1
X_14434_ _14502_/S vssd1 vssd1 vccd1 vccd1 _14443_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_156_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 io_dbus_rdata[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_4
X_17153_ _17204_/A vssd1 vssd1 vccd1 vccd1 _17167_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__15119__A2 _15116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput25 io_dbus_rdata[31] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_2
X_14365_ _14365_/A vssd1 vssd1 vccd1 vccd1 _18466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput36 io_ibus_inst[11] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10287__S1 _11113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11577_ _11598_/B _11476_/B _11366_/A vssd1 vssd1 vccd1 vccd1 _11599_/C sky130_fd_sc_hd__o21ba_1
XFILLER_156_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput47 io_ibus_inst[21] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__buf_2
Xinput58 io_ibus_inst[31] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_2
X_13316_ _13316_/A _13319_/B vssd1 vssd1 vccd1 vccd1 _13316_/X sky130_fd_sc_hd__or2_1
X_16104_ _16103_/X _19035_/Q _16113_/S vssd1 vssd1 vccd1 vccd1 _16105_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10061__B1 _09318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17084_ _16771_/X _19443_/Q _17086_/S vssd1 vssd1 vccd1 vccd1 _17085_/A sky130_fd_sc_hd__mux2_1
Xinput69 io_irq_m3_irq vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_6
X_10528_ _09927_/A _10518_/X _10527_/X _09307_/A _18436_/Q vssd1 vssd1 vccd1 vccd1
+ _12476_/B sky130_fd_sc_hd__a32o_4
XFILLER_170_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14296_ _14300_/A _14300_/B vssd1 vssd1 vccd1 vccd1 _14296_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13247_ _13185_/X _13245_/X _13246_/X _13232_/X vssd1 vssd1 vccd1 vccd1 _18359_/D
+ sky130_fd_sc_hd__o211a_1
X_16035_ _16116_/A vssd1 vssd1 vccd1 vccd1 _16135_/S sky130_fd_sc_hd__buf_8
X_10459_ _18438_/Q _09308_/A _09429_/A _10458_/X vssd1 vssd1 vccd1 vccd1 _12480_/A
+ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__14532__A _14565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13550__A1 _09106_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09626__A _18455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13178_ _13178_/A vssd1 vssd1 vccd1 vccd1 _13178_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13148__A _18620_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ _12129_/A vssd1 vssd1 vccd1 vccd1 _14178_/B sky130_fd_sc_hd__buf_2
XFILLER_69_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17986_ _18085_/A vssd1 vssd1 vccd1 vccd1 _18033_/A sky130_fd_sc_hd__buf_2
XFILLER_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13302__A1 _18282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19725_ _19725_/CLK _19725_/D vssd1 vssd1 vccd1 vccd1 _19725_/Q sky130_fd_sc_hd__dfxtp_1
X_16937_ _16937_/A vssd1 vssd1 vccd1 vccd1 _19377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17054__S _17058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10211__S1 _09978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19656_ _19723_/CLK _19656_/D vssd1 vssd1 vccd1 vccd1 _19656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16868_ _16868_/A vssd1 vssd1 vccd1 vccd1 _19347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18607_ _19329_/CLK _18607_/D vssd1 vssd1 vccd1 vccd1 _18607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15819_ _14761_/X _18917_/Q _15819_/S vssd1 vssd1 vccd1 vccd1 _15820_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19587_ _19587_/CLK _19587_/D vssd1 vssd1 vccd1 vccd1 _19587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16799_ _16799_/A vssd1 vssd1 vccd1 vccd1 _19323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09340_ _10387_/S vssd1 vssd1 vccd1 vccd1 _10277_/S sky130_fd_sc_hd__buf_4
X_18538_ _18548_/CLK _18538_/D vssd1 vssd1 vccd1 vccd1 _18538_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09904__S1 _09763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09271_ _10857_/B vssd1 vssd1 vccd1 vccd1 _11046_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_61_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18469_ _19080_/CLK _18469_/D vssd1 vssd1 vccd1 vccd1 _18469_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13369__A1 _18293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13369__B2 _18376_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16922__A _16990_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14318__B1 _14317_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15538__A _16793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09745__B1 _09414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15972__S _15972_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09271__A _10857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09607_ _09414_/A _09578_/Y _09581_/Y _09394_/A _09606_/X vssd1 vssd1 vccd1 vccd1
+ _09607_/X sky130_fd_sc_hd__o311a_2
XFILLER_44_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09538_ _09538_/A vssd1 vssd1 vccd1 vccd1 _09539_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10210__A _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09469_ _09463_/A _09466_/X _09468_/X _09459_/X vssd1 vssd1 vccd1 vccd1 _09469_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11500_ _11519_/A _11506_/A _11511_/C vssd1 vssd1 vccd1 vccd1 _13527_/B sky130_fd_sc_hd__or3_1
XFILLER_169_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12480_ _12480_/A _12483_/B vssd1 vssd1 vccd1 vccd1 _12480_/Y sky130_fd_sc_hd__nor2_1
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11431_ _18550_/Q vssd1 vssd1 vccd1 vccd1 _14582_/A sky130_fd_sc_hd__inv_2
XANTENNA__10269__S1 _09145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14150_ _14150_/A vssd1 vssd1 vccd1 vccd1 _14150_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11362_ _11362_/A _11375_/B vssd1 vssd1 vccd1 vccd1 _11478_/A sky130_fd_sc_hd__or2_1
XFILLER_165_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13101_ input69/X _13104_/B vssd1 vssd1 vccd1 vccd1 _13101_/X sky130_fd_sc_hd__or2_1
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10313_ _10313_/A _10313_/B vssd1 vssd1 vccd1 vccd1 _10313_/X sky130_fd_sc_hd__or2_1
X_14081_ _13821_/A _14073_/Y _14080_/Y vssd1 vssd1 vccd1 vccd1 _14081_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__16043__S _16049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11293_ _14875_/A vssd1 vssd1 vccd1 vccd1 _14737_/A sky130_fd_sc_hd__buf_2
X_13032_ _13033_/A _13033_/C _18323_/Q vssd1 vssd1 vccd1 vccd1 _13034_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_input52_A io_ibus_inst[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11695__B _13653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09446__A _09449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10244_ _10239_/X _10241_/Y _10243_/Y _10400_/A vssd1 vssd1 vccd1 vccd1 _10244_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10346__A1 _09430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16978__S _16986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09831__S0 _09928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17840_ _17840_/A vssd1 vssd1 vccd1 vccd1 _17849_/S sky130_fd_sc_hd__buf_4
XANTENNA__17663__A _17693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10441__S1 _10245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10175_ _10175_/A _10175_/B vssd1 vssd1 vccd1 vccd1 _10175_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15285__A1 _15162_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17771_ _15258_/X _17770_/Y _15263_/B vssd1 vssd1 vccd1 vccd1 _17771_/X sky130_fd_sc_hd__a21o_1
X_14983_ input16/X _14901_/X _14904_/X vssd1 vssd1 vccd1 vccd1 _14983_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_93_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19510_ _19659_/CLK _19510_/D vssd1 vssd1 vccd1 vccd1 _19510_/Q sky130_fd_sc_hd__dfxtp_1
X_16722_ _16722_/A vssd1 vssd1 vccd1 vccd1 _16735_/S sky130_fd_sc_hd__buf_4
X_13934_ _11751_/B _14319_/B _11460_/A vssd1 vssd1 vccd1 vccd1 _13934_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12600__A _12600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19441_ _19442_/CLK _19441_/D vssd1 vssd1 vccd1 vccd1 _19441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13415__B _18649_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16653_ _16653_/A vssd1 vssd1 vccd1 vccd1 _19278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13865_ _14278_/A vssd1 vssd1 vccd1 vccd1 _14314_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15604_ _15604_/A vssd1 vssd1 vccd1 vccd1 _18821_/D sky130_fd_sc_hd__clkbuf_1
X_12816_ _18254_/Q _12809_/C _12815_/Y vssd1 vssd1 vccd1 vccd1 _18254_/D sky130_fd_sc_hd__o21a_1
X_19372_ _19695_/CLK _19372_/D vssd1 vssd1 vccd1 vccd1 _19372_/Q sky130_fd_sc_hd__dfxtp_1
X_16584_ _16584_/A vssd1 vssd1 vccd1 vccd1 _19247_/D sky130_fd_sc_hd__clkbuf_1
X_13796_ _13796_/A vssd1 vssd1 vccd1 vccd1 _13797_/A sky130_fd_sc_hd__clkbuf_2
X_18323_ _19812_/CLK _18323_/D vssd1 vssd1 vccd1 vccd1 _18323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15535_ _16790_/A vssd1 vssd1 vccd1 vccd1 _15535_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12747_ _12791_/A _12751_/B _12747_/C vssd1 vssd1 vccd1 vccd1 _12748_/A sky130_fd_sc_hd__nor3_4
XANTENNA__17734__A0 _12757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16218__S _16224_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ _19872_/CLK _18254_/D vssd1 vssd1 vccd1 vccd1 _18254_/Q sky130_fd_sc_hd__dfxtp_1
X_12678_ _18349_/Q _15242_/A _12673_/X _12677_/X vssd1 vssd1 vccd1 vccd1 _12678_/X
+ sky130_fd_sc_hd__a211o_1
X_15466_ _18775_/Q _15210_/X _15470_/S vssd1 vssd1 vccd1 vccd1 _15467_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17205_ _18445_/Q _12634_/B _17218_/S vssd1 vssd1 vccd1 vccd1 _17205_/X sky130_fd_sc_hd__mux2_1
X_11629_ _14431_/B vssd1 vssd1 vccd1 vccd1 _11979_/A sky130_fd_sc_hd__clkbuf_2
X_14417_ _14417_/A vssd1 vssd1 vccd1 vccd1 _18484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18185_ _19849_/Q _18185_/B vssd1 vssd1 vccd1 vccd1 _18191_/C sky130_fd_sc_hd__and2_1
X_15397_ _15397_/A vssd1 vssd1 vccd1 vccd1 _15406_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__10034__B1 _10068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17136_ _11046_/A _13136_/X _17143_/S vssd1 vssd1 vccd1 vccd1 _17136_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09975__B1 _10107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14348_ _18461_/Q vssd1 vssd1 vccd1 vccd1 _17621_/A sky130_fd_sc_hd__buf_2
XFILLER_156_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17067_ _16743_/X _19435_/Q _17075_/S vssd1 vssd1 vccd1 vccd1 _17068_/A sky130_fd_sc_hd__mux2_1
X_14279_ _14278_/A _13959_/Y _14278_/Y _13737_/A vssd1 vssd1 vccd1 vccd1 _14279_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12326__A2 _14265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16018_ _16018_/A vssd1 vssd1 vccd1 vccd1 _16027_/S sky130_fd_sc_hd__buf_4
XFILLER_98_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15276__A1 _15149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14079__A2 _14074_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ _19774_/Q _17971_/C _17968_/Y vssd1 vssd1 vccd1 vccd1 _19774_/D sky130_fd_sc_hd__o21a_1
XFILLER_100_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19708_ _19708_/CLK _19708_/D vssd1 vssd1 vccd1 vccd1 _19708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19639_ _19639_/CLK _19639_/D vssd1 vssd1 vccd1 vccd1 _19639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17512__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15821__A _15878_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09889__S0 _09803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09323_ _10844_/A vssd1 vssd1 vccd1 vccd1 _10850_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10499__S1 _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09254_ _18529_/Q vssd1 vssd1 vccd1 vccd1 _09255_/A sky130_fd_sc_hd__inv_2
XFILLER_139_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09185_ _09712_/A vssd1 vssd1 vccd1 vccd1 _10210_/A sky130_fd_sc_hd__buf_2
XFILLER_119_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10576__A1 _10475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15268__A _15324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09813__S0 _09928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16798__S _16807_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10423__S1 _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_168_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11980_ _11980_/A vssd1 vssd1 vccd1 vccd1 _11980_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10931_ _09273_/A _10917_/X _10930_/X _11046_/B _18428_/Q vssd1 vssd1 vccd1 vccd1
+ _11070_/A sky130_fd_sc_hd__a32o_2
XFILLER_72_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17422__S _17424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13650_ _13650_/A vssd1 vssd1 vccd1 vccd1 _13993_/A sky130_fd_sc_hd__clkbuf_1
X_10862_ _19248_/Q _19019_/Q _18950_/Q _19344_/Q _10614_/X _10616_/X vssd1 vssd1 vccd1
+ vccd1 _10863_/B sky130_fd_sc_hd__mux4_2
XFILLER_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _13415_/A _18637_/Q vssd1 vssd1 vccd1 vccd1 _12601_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12253__A1 _12246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16519__A1 _15510_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13581_ _13712_/B vssd1 vssd1 vccd1 vccd1 _13785_/A sky130_fd_sc_hd__buf_2
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10875__A _10875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10793_ _10793_/A vssd1 vssd1 vccd1 vccd1 _10793_/X sky130_fd_sc_hd__clkbuf_2
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15320_ _18712_/Q _15213_/X _15322_/S vssd1 vssd1 vccd1 vccd1 _15321_/A sky130_fd_sc_hd__mux2_1
X_12532_ _12532_/A vssd1 vssd1 vccd1 vccd1 _12643_/A sky130_fd_sc_hd__clkbuf_2
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15251_ _11759_/B _13149_/X _17143_/S vssd1 vssd1 vccd1 vccd1 _15251_/X sky130_fd_sc_hd__mux2_1
X_12463_ _12463_/A _12466_/B vssd1 vssd1 vccd1 vccd1 _12464_/A sky130_fd_sc_hd__and2_1
X_11414_ _11423_/A _12519_/A _12791_/B vssd1 vssd1 vccd1 vccd1 _12563_/A sky130_fd_sc_hd__nor3_1
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14202_ _13927_/X _14199_/Y _14201_/X _13982_/X vssd1 vssd1 vccd1 vccd1 _14202_/X
+ sky130_fd_sc_hd__a211o_1
X_15182_ _18664_/Q _15181_/X _15185_/S vssd1 vssd1 vccd1 vccd1 _15183_/A sky130_fd_sc_hd__mux2_1
X_12394_ _11790_/A _12392_/Y _12414_/B _12116_/A vssd1 vssd1 vccd1 vccd1 _12394_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_137_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10567__A1 _09454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14133_ _12041_/Y _14070_/X _14132_/X _14099_/X vssd1 vssd1 vccd1 vccd1 _14133_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__15178__A _16680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11345_ _11374_/A _11375_/A _11519_/B vssd1 vssd1 vccd1 vccd1 _11345_/Y sky130_fd_sc_hd__nor3_1
XFILLER_4_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10814__S _11028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18941_ _19724_/CLK _18941_/D vssd1 vssd1 vccd1 vccd1 _18941_/Q sky130_fd_sc_hd__dfxtp_1
X_14064_ _13970_/S _13953_/X _13899_/X vssd1 vssd1 vccd1 vccd1 _14220_/B sky130_fd_sc_hd__o21ai_1
X_11276_ _11149_/A _11225_/X _11151_/A vssd1 vssd1 vccd1 vccd1 _11276_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_140_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13015_ _13015_/A _18317_/Q _13015_/C vssd1 vssd1 vccd1 vccd1 _13016_/C sky130_fd_sc_hd__and3_1
XFILLER_79_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17393__A _17461_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10227_ _10227_/A vssd1 vssd1 vccd1 vccd1 _11119_/A sky130_fd_sc_hd__buf_2
X_18872_ _19331_/CLK _18872_/D vssd1 vssd1 vccd1 vccd1 _18872_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10115__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16501__S _16501_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17823_ _15194_/X _19713_/Q _17827_/S vssd1 vssd1 vccd1 vccd1 _17824_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10158_ _18771_/Q _19000_/Q _18931_/Q _19229_/Q _10256_/S _09145_/A vssd1 vssd1 vccd1
+ vccd1 _10159_/B sky130_fd_sc_hd__mux4_1
XFILLER_121_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17754_ _17730_/X _13387_/X _17724_/X vssd1 vssd1 vccd1 vccd1 _17754_/X sky130_fd_sc_hd__a21bo_1
X_14966_ _14966_/A vssd1 vssd1 vccd1 vccd1 _18607_/D sky130_fd_sc_hd__clkbuf_1
X_10089_ _10120_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10089_/X sky130_fd_sc_hd__or2_1
XFILLER_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10178__S0 _09721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16705_ _16705_/A vssd1 vssd1 vccd1 vccd1 _16705_/X sky130_fd_sc_hd__clkbuf_2
X_13917_ _13916_/X _13897_/X _14121_/S vssd1 vssd1 vccd1 vccd1 _13917_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17685_ _17691_/B _17685_/B vssd1 vssd1 vccd1 vccd1 _17685_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16737__A _16737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14897_ _18442_/Q _12554_/B _14981_/S vssd1 vssd1 vccd1 vccd1 _14897_/X sky130_fd_sc_hd__mux2_1
X_19424_ _19717_/CLK _19424_/D vssd1 vssd1 vccd1 vccd1 _19424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16636_ _16636_/A vssd1 vssd1 vccd1 vccd1 _19273_/D sky130_fd_sc_hd__clkbuf_1
X_13848_ _13848_/A vssd1 vssd1 vccd1 vccd1 _13848_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19355_ _19613_/CLK _19355_/D vssd1 vssd1 vccd1 vccd1 _19355_/Q sky130_fd_sc_hd__dfxtp_1
X_16567_ _19239_/Q _15580_/X _16569_/S vssd1 vssd1 vccd1 vccd1 _16568_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10785__A _10785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13779_ _13838_/A vssd1 vssd1 vccd1 vccd1 _14121_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18306_ _18329_/CLK _18306_/D vssd1 vssd1 vccd1 vccd1 _18306_/Q sky130_fd_sc_hd__dfxtp_1
X_15518_ _15518_/A vssd1 vssd1 vccd1 vccd1 _18793_/D sky130_fd_sc_hd__clkbuf_1
X_19286_ _19414_/CLK _19286_/D vssd1 vssd1 vccd1 vccd1 _19286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16498_ _16498_/A vssd1 vssd1 vccd1 vccd1 _19208_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15787__S _15791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18237_ _18239_/B _18239_/C _18170_/X vssd1 vssd1 vccd1 vccd1 _18237_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_90_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15449_ _15449_/A vssd1 vssd1 vccd1 vccd1 _18767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18168_ _18197_/A _18175_/C vssd1 vssd1 vccd1 vccd1 _18168_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11755__B1 _17221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17119_ _16822_/X _19459_/Q _17119_/S vssd1 vssd1 vccd1 vccd1 _17120_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18099_ _19819_/Q _18096_/B _18098_/Y vssd1 vssd1 vccd1 vccd1 _19819_/D sky130_fd_sc_hd__o21a_1
XFILLER_143_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12505__A _12505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10653__S1 _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09941_ _19524_/Q _19138_/Q _19588_/Q _18744_/Q _09866_/X _09881_/X vssd1 vssd1 vccd1
+ vccd1 _09942_/B sky130_fd_sc_hd__mux4_1
XFILLER_143_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17507__S _17507_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16411__S _16413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09872_ _18874_/Q _19332_/Q _09872_/S vssd1 vssd1 vccd1 vccd1 _09873_/A sky130_fd_sc_hd__mux2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14720__A _16744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09814__A _09814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17242__S _17245_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09306_ _09306_/A vssd1 vssd1 vccd1 vccd1 _09307_/A sky130_fd_sc_hd__buf_2
XFILLER_167_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17174__A1 _13259_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09237_ _09237_/A _09237_/B vssd1 vssd1 vccd1 vccd1 _09237_/X sky130_fd_sc_hd__or2_1
XFILLER_155_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_94_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16382__A _16428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13735__A1 _11046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09168_ _09168_/A vssd1 vssd1 vccd1 vccd1 _09169_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_107_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10644__S1 _10634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09099_ _18558_/Q vssd1 vssd1 vccd1 vccd1 _11321_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_150_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11130_ _11130_/A _12481_/A vssd1 vssd1 vccd1 vccd1 _11130_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14160__A1 _12096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061_ _19629_/Q _19046_/Q _19083_/Q _18689_/Q _10710_/A _09480_/A vssd1 vssd1 vccd1
+ vccd1 _11062_/B sky130_fd_sc_hd__mux4_2
XFILLER_1_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16321__S _16329_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10012_ _10115_/A _10011_/X _10093_/A vssd1 vssd1 vccd1 vccd1 _10012_/X sky130_fd_sc_hd__a21o_1
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14820_ _16670_/A vssd1 vssd1 vccd1 vccd1 _16774_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input15_A io_dbus_rdata[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14751_ input26/X _14703_/X _14750_/Y _14711_/X vssd1 vssd1 vccd1 vccd1 _16651_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11963_ _12020_/C vssd1 vssd1 vccd1 vccd1 _11963_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13702_ _13702_/A _13996_/B vssd1 vssd1 vccd1 vccd1 _13703_/A sky130_fd_sc_hd__nand2_1
X_17470_ _19599_/Q _16648_/X _17474_/S vssd1 vssd1 vccd1 vccd1 _17471_/A sky130_fd_sc_hd__mux2_1
X_10914_ _18755_/Q _18984_/Q _18915_/Q _19213_/Q _10959_/A _10910_/A vssd1 vssd1 vccd1
+ vccd1 _10915_/B sky130_fd_sc_hd__mux4_1
X_14682_ _14694_/A _14682_/B vssd1 vssd1 vccd1 vccd1 _14683_/A sky130_fd_sc_hd__and2_1
XFILLER_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11894_ _12057_/A _14026_/A _11867_/B vssd1 vssd1 vccd1 vccd1 _11895_/B sky130_fd_sc_hd__a21oi_2
X_16421_ _16421_/A vssd1 vssd1 vccd1 vccd1 _19174_/D sky130_fd_sc_hd__clkbuf_1
X_13633_ _11784_/A _12372_/A _13659_/S vssd1 vssd1 vccd1 vccd1 _13633_/X sky130_fd_sc_hd__mux2_1
X_10845_ _10899_/A _10842_/X _10844_/X _10793_/X vssd1 vssd1 vccd1 vccd1 _10846_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19140_ _19657_/CLK _19140_/D vssd1 vssd1 vccd1 vccd1 _19140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16352_ _16352_/A vssd1 vssd1 vccd1 vccd1 _19144_/D sky130_fd_sc_hd__clkbuf_1
X_10776_ _19409_/Q _19185_/Q _19702_/Q _19153_/Q _10724_/X _10713_/X vssd1 vssd1 vccd1
+ vccd1 _10776_/X sky130_fd_sc_hd__mux4_1
X_13564_ _13564_/A vssd1 vssd1 vccd1 vccd1 _18425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10332__S0 _10328_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15303_ _18704_/Q _15187_/X _15311_/S vssd1 vssd1 vccd1 vccd1 _15304_/A sky130_fd_sc_hd__mux2_1
X_19071_ _19721_/CLK _19071_/D vssd1 vssd1 vccd1 vccd1 _19071_/Q sky130_fd_sc_hd__dfxtp_1
X_12515_ _19808_/Q vssd1 vssd1 vccd1 vccd1 _18067_/B sky130_fd_sc_hd__clkbuf_2
X_13495_ _18406_/Q _12757_/X _13497_/S vssd1 vssd1 vccd1 vccd1 _13496_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16283_ _16134_/X _19114_/Q _16283_/S vssd1 vssd1 vccd1 vccd1 _16284_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18022_ _18023_/A _18023_/B _18021_/Y vssd1 vssd1 vccd1 vccd1 _19793_/D sky130_fd_sc_hd__o21a_1
XANTENNA__15400__S _15406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12446_ _14332_/B _12446_/B vssd1 vssd1 vccd1 vccd1 _12447_/B sky130_fd_sc_hd__or2_1
X_15234_ _15234_/A vssd1 vssd1 vccd1 vccd1 _18680_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15165_ _16667_/A vssd1 vssd1 vccd1 vccd1 _15165_/X sky130_fd_sc_hd__clkbuf_2
X_12377_ _12419_/A _12377_/B vssd1 vssd1 vccd1 vccd1 _14300_/A sky130_fd_sc_hd__nand2_2
XFILLER_126_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10635__S1 _10634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14116_ _13726_/X _14105_/Y _14114_/X _14115_/X vssd1 vssd1 vccd1 vccd1 _14116_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA_output83_A _12163_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11328_ _11513_/A _11514_/A _18581_/Q _18584_/Q vssd1 vssd1 vccd1 vccd1 _11640_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_140_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15096_ _15125_/A vssd1 vssd1 vccd1 vccd1 _15111_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_153_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18924_ _19707_/CLK _18924_/D vssd1 vssd1 vccd1 vccd1 _18924_/Q sky130_fd_sc_hd__dfxtp_1
X_14047_ _14042_/Y _14044_/Y _14046_/X vssd1 vssd1 vccd1 vccd1 _14047_/X sky130_fd_sc_hd__a21o_1
X_11259_ _11080_/C _11248_/Y _11250_/Y _11255_/X _11258_/X vssd1 vssd1 vccd1 vccd1
+ _11261_/C sky130_fd_sc_hd__a2111o_1
XANTENNA__14540__A _15339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10399__S0 _10277_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18855_ _19539_/CLK _18855_/D vssd1 vssd1 vccd1 vccd1 _18855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17806_ _17806_/A vssd1 vssd1 vccd1 vccd1 _19705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18786_ _19534_/CLK _18786_/D vssd1 vssd1 vccd1 vccd1 _18786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15998_ _15998_/A vssd1 vssd1 vccd1 vccd1 _18997_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13111__C1 _13102_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17737_ _17737_/A _18482_/Q _17737_/C vssd1 vssd1 vccd1 vccd1 _17743_/B sky130_fd_sc_hd__or3_1
XANTENNA__13662__A0 _12355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_161_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19691_/CLK sky130_fd_sc_hd__clkbuf_16
X_14949_ _14811_/X _14945_/X _14947_/X _14948_/X vssd1 vssd1 vccd1 vccd1 _16705_/A
+ sky130_fd_sc_hd__o31a_2
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17062__S _17062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17668_ _17662_/A _17667_/C _14861_/A vssd1 vssd1 vccd1 vccd1 _17669_/B sky130_fd_sc_hd__o21ai_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10571__S0 _11088_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19407_ _19700_/CLK _19407_/D vssd1 vssd1 vccd1 vccd1 _19407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16619_ _19265_/Q vssd1 vssd1 vccd1 vccd1 _16620_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_126_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17599_ _19657_/Q _16835_/A _17601_/S vssd1 vssd1 vccd1 vccd1 _17600_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19338_ _19648_/CLK _19338_/D vssd1 vssd1 vccd1 vccd1 _19338_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_176_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19702_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19269_ _19622_/CLK _19269_/D vssd1 vssd1 vccd1 vccd1 _19269_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10874__S1 _10616_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14715__A _18533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09809__A _09872_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10626__S1 _10548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_114_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19733_/CLK sky130_fd_sc_hd__clkbuf_16
X_09924_ _09624_/A _09624_/B _09425_/Y vssd1 vssd1 vccd1 vccd1 _09925_/A sky130_fd_sc_hd__a21oi_1
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09544__A _09793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ _19526_/Q _19140_/Q _19590_/Q _18746_/Q _09163_/A _09843_/A vssd1 vssd1 vccd1
+ vccd1 _09856_/B sky130_fd_sc_hd__mux4_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A io_dbus_rdata[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11900__B1 _19737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09786_ _09217_/A _09776_/X _09778_/X _09785_/X _09854_/A vssd1 vssd1 vccd1 vccd1
+ _09786_/X sky130_fd_sc_hd__a221o_4
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_129_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _18487_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10467__B1 _09454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _09274_/A _10620_/X _10629_/X _09281_/A _18434_/Q vssd1 vssd1 vccd1 vccd1
+ _11077_/A sky130_fd_sc_hd__a32o_2
XFILLER_41_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10561_ _09170_/A _10560_/X _09451_/A vssd1 vssd1 vccd1 vccd1 _10561_/X sky130_fd_sc_hd__a21o_1
XFILLER_155_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10865__S1 _10740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16316__S _16318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12300_ _12298_/Y _12299_/X _17886_/A vssd1 vssd1 vccd1 vccd1 _12300_/X sky130_fd_sc_hd__o21a_1
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13280_ _18363_/Q _13295_/B vssd1 vssd1 vccd1 vccd1 _13280_/X sky130_fd_sc_hd__or2_1
X_10492_ _10591_/A _10492_/B vssd1 vssd1 vccd1 vccd1 _10492_/X sky130_fd_sc_hd__or2_1
X_12231_ _18512_/Q _12259_/B _12259_/C vssd1 vssd1 vccd1 vccd1 _12231_/X sky130_fd_sc_hd__or3_1
XANTENNA__13184__A2 _13182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14381__A1 _18504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10617__S1 _10616_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11195__A1 _09317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12162_ _12141_/A _12141_/B _12138_/A vssd1 vssd1 vccd1 vccd1 _12163_/B sky130_fd_sc_hd__a21oi_2
XFILLER_122_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11984__A _11984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ _11113_/A _11113_/B vssd1 vssd1 vccd1 vccd1 _11113_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14133__A1 _12041_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16970_ _16970_/A vssd1 vssd1 vccd1 vccd1 _19392_/D sky130_fd_sc_hd__clkbuf_1
X_12093_ _19740_/Q _19741_/Q _19742_/Q _12093_/D vssd1 vssd1 vccd1 vccd1 _12094_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_122_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11044_ _11037_/Y _11039_/Y _11041_/Y _11043_/Y _19695_/Q vssd1 vssd1 vccd1 vccd1
+ _11044_/X sky130_fd_sc_hd__o221a_2
XANTENNA__09454__A _09454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15921_ _15921_/A vssd1 vssd1 vccd1 vccd1 _18962_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11042__S1 _10920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16986__S _16986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18640_ _19804_/CLK _18640_/D vssd1 vssd1 vccd1 vccd1 _18640_/Q sky130_fd_sc_hd__dfxtp_1
X_15852_ _14940_/X _18932_/Q _15852_/S vssd1 vssd1 vccd1 vccd1 _15853_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14803_ _14842_/A _14803_/B vssd1 vssd1 vccd1 vccd1 _14804_/A sky130_fd_sc_hd__or2_2
XFILLER_91_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13644__A0 _12510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18571_ _18578_/CLK _18571_/D vssd1 vssd1 vccd1 vccd1 _18571_/Q sky130_fd_sc_hd__dfxtp_1
X_15783_ _14951_/X _18901_/Q _15791_/S vssd1 vssd1 vccd1 vccd1 _15784_/A sky130_fd_sc_hd__mux2_1
X_12995_ _18310_/Q _18312_/Q _18311_/Q _12995_/D vssd1 vssd1 vccd1 vccd1 _13006_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16287__A _16355_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17522_ _17522_/A vssd1 vssd1 vccd1 vccd1 _19622_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15191__A _16693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14734_ _14873_/A vssd1 vssd1 vccd1 vccd1 _14958_/A sky130_fd_sc_hd__clkbuf_2
X_11946_ _12030_/B vssd1 vssd1 vccd1 vccd1 _14075_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_93_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19859_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14519__B _14519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17453_ _16832_/X _19592_/Q _17457_/S vssd1 vssd1 vccd1 vccd1 _17454_/A sky130_fd_sc_hd__mux2_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ _14566_/A _12660_/A _14640_/A input47/X vssd1 vssd1 vccd1 vccd1 _15954_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _11844_/B _11874_/Y _11846_/A _11876_/X vssd1 vssd1 vccd1 vccd1 _11877_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_32_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16404_ _16415_/A vssd1 vssd1 vccd1 vccd1 _16413_/S sky130_fd_sc_hd__buf_6
X_13616_ _14045_/B _13615_/Y _13681_/S vssd1 vssd1 vccd1 vccd1 _13616_/X sky130_fd_sc_hd__mux2_1
X_17384_ _17384_/A vssd1 vssd1 vccd1 vccd1 _19561_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10828_ _10830_/A _10826_/X _10827_/X vssd1 vssd1 vccd1 vccd1 _10828_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11958__A0 _11956_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14596_ _14612_/A _14596_/B vssd1 vssd1 vccd1 vccd1 _18554_/D sky130_fd_sc_hd__nand2_1
X_19123_ _19638_/CLK _19123_/D vssd1 vssd1 vccd1 vccd1 _19123_/Q sky130_fd_sc_hd__dfxtp_1
X_16335_ _16335_/A vssd1 vssd1 vccd1 vccd1 _19136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13547_ _16212_/C _13537_/X _13546_/X vssd1 vssd1 vccd1 vccd1 _13548_/B sky130_fd_sc_hd__a21bo_1
X_10759_ _19603_/Q _19441_/Q _18887_/Q _18657_/Q _10836_/A _09353_/A vssd1 vssd1 vccd1
+ vccd1 _10760_/B sky130_fd_sc_hd__mux4_1
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18007__A _18033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09629__A _09629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19054_ _19635_/CLK _19054_/D vssd1 vssd1 vccd1 vccd1 _19054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16266_ _16109_/X _19106_/Q _16268_/S vssd1 vssd1 vccd1 vccd1 _16267_/A sky130_fd_sc_hd__mux2_1
X_13478_ _18398_/Q _13307_/X _13486_/S vssd1 vssd1 vccd1 vccd1 _13479_/A sky130_fd_sc_hd__mux2_1
X_18005_ _19786_/Q _18006_/C hold2/A vssd1 vssd1 vccd1 vccd1 _18007_/B sky130_fd_sc_hd__a21oi_1
X_15217_ _18675_/Q _15216_/X _15217_/S vssd1 vssd1 vccd1 vccd1 _15218_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12429_ _12385_/A _12385_/B _12404_/B _12384_/A vssd1 vssd1 vccd1 vccd1 _12430_/B
+ sky130_fd_sc_hd__a211o_1
X_16197_ _16115_/X _19071_/Q _16205_/S vssd1 vssd1 vccd1 vccd1 _16198_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_31_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19326_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15148_ _15148_/A vssd1 vssd1 vccd1 vccd1 _18653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15079_ _15079_/A vssd1 vssd1 vccd1 vccd1 _15092_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__12135__A0 _10196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09364__A _09364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18907_ _19722_/CLK _18907_/D vssd1 vssd1 vccd1 vccd1 _18907_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16896__S _16902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_46_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19554_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_42_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17581__A _17592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09640_ _09640_/A _09640_/B vssd1 vssd1 vccd1 vccd1 _09640_/X sky130_fd_sc_hd__or2_1
XFILLER_83_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18838_ _19003_/CLK _18838_/D vssd1 vssd1 vccd1 vccd1 _18838_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10303__A _10309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09571_ _09649_/A _09571_/B vssd1 vssd1 vccd1 vccd1 _09571_/X sky130_fd_sc_hd__or2_1
X_18769_ _19581_/CLK _18769_/D vssd1 vssd1 vccd1 vccd1 _18769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15305__S _15311_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13614__A _13614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10847__S1 _10634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11788__B _11788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14164__B _14168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15975__S _15983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13323__C1 _13317_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09907_ _18840_/Q _19394_/Q _19556_/Q _18808_/Q _09976_/A _09783_/A vssd1 vssd1 vccd1
+ vccd1 _09908_/B sky130_fd_sc_hd__mux4_1
XFILLER_99_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13874__B1 _13873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09838_ _18450_/Q vssd1 vssd1 vccd1 vccd1 _09838_/Y sky130_fd_sc_hd__inv_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09769_ _09769_/A vssd1 vssd1 vccd1 vccd1 _09783_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11800_ _11827_/B _11798_/Y _11799_/X _15262_/A vssd1 vssd1 vccd1 vccd1 _11800_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _12765_/X _12779_/X _12780_/S vssd1 vssd1 vccd1 vccd1 _12780_/X sky130_fd_sc_hd__mux2_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _19731_/Q _11705_/X _11713_/X _11730_/X vssd1 vssd1 vccd1 vccd1 _17860_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _18497_/Q _19735_/Q _14454_/S vssd1 vssd1 vccd1 vccd1 _14451_/A sky130_fd_sc_hd__mux2_1
X_11662_ _19730_/Q _13529_/A vssd1 vssd1 vccd1 vccd1 _11752_/C sky130_fd_sc_hd__and2_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _14514_/A vssd1 vssd1 vccd1 vccd1 _13401_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_168_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10613_ _10992_/A vssd1 vssd1 vccd1 vccd1 _10873_/A sky130_fd_sc_hd__buf_2
XFILLER_168_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16046__S _16049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11593_ _11593_/A vssd1 vssd1 vccd1 vccd1 _12259_/C sky130_fd_sc_hd__clkbuf_2
X_14381_ _17683_/A _18504_/Q _14381_/S vssd1 vssd1 vccd1 vccd1 _14382_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16120_ _16119_/X _19040_/Q _16129_/S vssd1 vssd1 vccd1 vccd1 _16121_/A sky130_fd_sc_hd__mux2_1
X_13332_ _19845_/Q _12736_/X _13331_/X vssd1 vssd1 vccd1 vccd1 _14958_/D sky130_fd_sc_hd__a21o_1
X_10544_ _19413_/Q _19189_/Q _19706_/Q _19157_/Q _10558_/S _10367_/A vssd1 vssd1 vccd1
+ vccd1 _10544_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09449__A _09449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11698__B _13667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14074__B _14074_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15885__S _15891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16051_ _16761_/A vssd1 vssd1 vccd1 vccd1 _16051_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13263_ _18361_/Q _13295_/B vssd1 vssd1 vccd1 vccd1 _13263_/X sky130_fd_sc_hd__or2_1
X_10475_ _10475_/A _10475_/B vssd1 vssd1 vccd1 vccd1 _10475_/X sky130_fd_sc_hd__or2_1
XFILLER_108_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15002_ _18482_/Q _18483_/Q _15002_/C vssd1 vssd1 vccd1 vccd1 _15015_/B sky130_fd_sc_hd__and3_1
X_12214_ _19680_/Q vssd1 vssd1 vccd1 vccd1 _12214_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13194_ _18308_/Q _13178_/A _12664_/A _19797_/Q _13193_/X vssd1 vssd1 vccd1 vccd1
+ _13194_/X sky130_fd_sc_hd__a221o_1
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19810_ _19810_/CLK _19810_/D vssd1 vssd1 vccd1 vccd1 _19810_/Q sky130_fd_sc_hd__dfxtp_1
X_12145_ _12145_/A _12215_/C vssd1 vssd1 vccd1 vccd1 _12145_/X sky130_fd_sc_hd__or2_1
XANTENNA__12603__A _12603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14657__A2 _12660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09184__A _09184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12076_ _12091_/A _12074_/Y _12123_/C _11859_/X vssd1 vssd1 vccd1 vccd1 _12076_/Y
+ sky130_fd_sc_hd__o31ai_1
X_19741_ _19753_/CLK _19741_/D vssd1 vssd1 vccd1 vccd1 _19741_/Q sky130_fd_sc_hd__dfxtp_1
X_16953_ _16790_/X _19385_/Q _16953_/S vssd1 vssd1 vccd1 vccd1 _16954_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15904_ _15950_/S vssd1 vssd1 vccd1 vccd1 _15913_/S sky130_fd_sc_hd__buf_2
X_11027_ _18586_/Q _19275_/Q _11027_/S vssd1 vssd1 vccd1 vccd1 _11027_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17605__S _17605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19672_ _19687_/CLK _19672_/D vssd1 vssd1 vccd1 vccd1 _19672_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_38_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09533__B2 _09532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16884_ _16884_/A vssd1 vssd1 vccd1 vccd1 _19354_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15606__A1 _15506_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18623_ _18623_/CLK _18623_/D vssd1 vssd1 vccd1 vccd1 _18623_/Q sky130_fd_sc_hd__dfxtp_2
X_15835_ _14847_/X _18924_/Q _15841_/S vssd1 vssd1 vccd1 vccd1 _15836_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18554_ _19733_/CLK _18554_/D vssd1 vssd1 vccd1 vccd1 _18554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15766_ _15766_/A vssd1 vssd1 vccd1 vccd1 _18893_/D sky130_fd_sc_hd__clkbuf_1
X_12978_ _18307_/Q vssd1 vssd1 vccd1 vccd1 _12982_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _19615_/Q _16699_/X _17507_/S vssd1 vssd1 vccd1 vccd1 _17506_/A sky130_fd_sc_hd__mux2_1
X_14717_ _16919_/A _16919_/B _15134_/A vssd1 vssd1 vccd1 vccd1 _16744_/A sky130_fd_sc_hd__or3b_4
XFILLER_61_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11929_ _12016_/S vssd1 vssd1 vccd1 vccd1 _12408_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18485_ _19686_/CLK _18485_/D vssd1 vssd1 vccd1 vccd1 _18485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15697_ _18863_/Q _15535_/X _15697_/S vssd1 vssd1 vccd1 vccd1 _15698_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17436_ _17436_/A vssd1 vssd1 vccd1 vccd1 _19584_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14648_ _14648_/A vssd1 vssd1 vccd1 vccd1 _14648_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11889__A _17221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ _17367_/A vssd1 vssd1 vccd1 vccd1 _19553_/D sky130_fd_sc_hd__clkbuf_1
X_14579_ _18548_/Q _14577_/X _14578_/X _14573_/X vssd1 vssd1 vccd1 vccd1 _18548_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14265__A _14265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10793__A _10793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10829__S1 _10813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19106_ _19718_/CLK _19106_/D vssd1 vssd1 vccd1 vccd1 _19106_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09359__A _11189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16318_ _16080_/X _19129_/Q _16318_/S vssd1 vssd1 vccd1 vccd1 _16319_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11800__C1 _15262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17298_ _19523_/Q _16712_/X _17302_/S vssd1 vssd1 vccd1 vccd1 _17299_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19037_ _19427_/CLK _19037_/D vssd1 vssd1 vccd1 vccd1 _19037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16249_ _16083_/X _19098_/Q _16257_/S vssd1 vssd1 vccd1 vccd1 _16250_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11159__A1 _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput102 _11846_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[7] sky130_fd_sc_hd__buf_2
Xoutput113 _12479_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[11] sky130_fd_sc_hd__buf_2
XFILLER_127_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput124 _12492_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[21] sky130_fd_sc_hd__buf_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15808__B _16503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput135 _12505_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[31] sky130_fd_sc_hd__buf_2
XFILLER_99_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput146 _17876_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[11] sky130_fd_sc_hd__buf_2
XFILLER_82_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput157 _12225_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[21] sky130_fd_sc_hd__buf_2
XANTENNA__15096__A _15125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput168 _12457_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[31] sky130_fd_sc_hd__buf_2
XFILLER_99_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12513__A _12766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09094__A _09094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14431__C _14431_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11006__S1 _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11129__A _11130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10765__S0 _10650_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09623_ _09612_/Y _09617_/Y _09619_/Y _09622_/Y _09403_/A vssd1 vssd1 vccd1 vccd1
+ _09623_/X sky130_fd_sc_hd__o221a_2
XFILLER_37_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09554_ _09554_/A vssd1 vssd1 vccd1 vccd1 _09642_/A sky130_fd_sc_hd__buf_2
XFILLER_83_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09485_ _10392_/A _09485_/B vssd1 vssd1 vccd1 vccd1 _09485_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17250__S _17258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15533__A0 _18798_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10260_ _19419_/Q _19195_/Q _19712_/Q _19163_/Q _09794_/A _09697_/A vssd1 vssd1 vccd1
+ vccd1 _10260_/X sky130_fd_sc_hd__mux4_2
XFILLER_152_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10191_ _10177_/A _10188_/X _10190_/X vssd1 vssd1 vccd1 vccd1 _10191_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13950_ _13950_/A vssd1 vssd1 vccd1 vccd1 _13950_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12901_ _12910_/D _12897_/B _12900_/Y vssd1 vssd1 vccd1 vccd1 _18279_/D sky130_fd_sc_hd__o21a_1
XANTENNA__11981__B _19737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13881_ _13879_/X _13993_/B _13881_/S vssd1 vssd1 vccd1 vccd1 _13881_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15620_ _15620_/A vssd1 vssd1 vccd1 vccd1 _18828_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _18260_/Q _18259_/Q _18258_/Q _12832_/D vssd1 vssd1 vccd1 vccd1 _12842_/D
+ sky130_fd_sc_hd__and4_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10508__S0 _10387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _16806_/A vssd1 vssd1 vccd1 vccd1 _15551_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _14519_/B vssd1 vssd1 vccd1 vccd1 _12763_/X sky130_fd_sc_hd__buf_2
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17210__A0 _19489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11181__S0 _10185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _18521_/Q _19759_/Q _14502_/S vssd1 vssd1 vccd1 vccd1 _14503_/A sky130_fd_sc_hd__mux2_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _19472_/CLK _18270_/D vssd1 vssd1 vccd1 vccd1 _18270_/Q sky130_fd_sc_hd__dfxtp_1
X_11714_ _17611_/B vssd1 vssd1 vccd1 vccd1 _15262_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _15482_/A vssd1 vssd1 vccd1 vccd1 _18782_/D sky130_fd_sc_hd__clkbuf_1
X_12694_ _13042_/A vssd1 vssd1 vccd1 vccd1 _17882_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17221_ _17221_/A vssd1 vssd1 vccd1 vccd1 _17235_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13378__A2 _13376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14433_ _14591_/B vssd1 vssd1 vccd1 vccd1 _14502_/S sky130_fd_sc_hd__buf_2
X_11645_ _13584_/C _11645_/B _13584_/D _13571_/C vssd1 vssd1 vccd1 vccd1 _12005_/A
+ sky130_fd_sc_hd__nor4b_4
XFILLER_52_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17152_ _17152_/A vssd1 vssd1 vccd1 vccd1 _19472_/D sky130_fd_sc_hd__clkbuf_1
X_14364_ _17645_/A _18498_/Q _14367_/S vssd1 vssd1 vccd1 vccd1 _14365_/A sky130_fd_sc_hd__mux2_1
Xinput15 io_dbus_rdata[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_2
XFILLER_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput26 io_dbus_rdata[3] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11576_ _11497_/A _11575_/Y _15079_/A _11556_/A vssd1 vssd1 vccd1 vccd1 _11576_/X
+ sky130_fd_sc_hd__a2bb2o_1
Xinput37 io_ibus_inst[12] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10597__C1 _09314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput48 io_ibus_inst[22] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_4
X_16103_ _16813_/A vssd1 vssd1 vccd1 vccd1 _16103_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13315_ _12598_/B _13311_/X _13314_/X _13282_/X vssd1 vssd1 vccd1 vccd1 _18367_/D
+ sky130_fd_sc_hd__o211a_1
Xinput59 io_ibus_inst[3] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_1
X_17083_ _17083_/A vssd1 vssd1 vccd1 vccd1 _19442_/D sky130_fd_sc_hd__clkbuf_1
X_10527_ _10520_/X _10522_/X _10524_/X _10526_/X _09392_/A vssd1 vssd1 vccd1 vccd1
+ _10527_/X sky130_fd_sc_hd__a221o_2
X_14295_ _18453_/Q _11460_/A _14284_/Y _14294_/X vssd1 vssd1 vccd1 vccd1 _18453_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_171_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16034_ _16847_/A _17064_/B vssd1 vssd1 vccd1 vccd1 _16116_/A sky130_fd_sc_hd__or2_2
X_13246_ _13246_/A _13246_/B vssd1 vssd1 vccd1 vccd1 _13246_/X sky130_fd_sc_hd__or2_1
XFILLER_6_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10458_ _09402_/A _10445_/X _10457_/X vssd1 vssd1 vccd1 vccd1 _10458_/X sky130_fd_sc_hd__a21o_2
XFILLER_171_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13177_ _19860_/Q _12604_/X _12749_/A _18031_/B vssd1 vssd1 vccd1 vccd1 _13177_/X
+ sky130_fd_sc_hd__a22o_1
X_10389_ _18600_/Q _19289_/Q _10389_/S vssd1 vssd1 vccd1 vccd1 _10390_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10995__S0 _10959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13148__B _13148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ _12155_/A _12128_/B vssd1 vssd1 vccd1 vccd1 _12129_/A sky130_fd_sc_hd__nand2_1
X_17985_ _19780_/Q _17988_/C _17984_/Y vssd1 vssd1 vccd1 vccd1 _19780_/D sky130_fd_sc_hd__o21a_1
XFILLER_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19724_ _19724_/CLK _19724_/D vssd1 vssd1 vccd1 vccd1 _19724_/Q sky130_fd_sc_hd__dfxtp_1
X_16936_ _16765_/X _19377_/Q _16942_/S vssd1 vssd1 vccd1 vccd1 _16937_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12059_ _14140_/B _12059_/B vssd1 vssd1 vccd1 vccd1 _12063_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__18020__A _18207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09642__A _09642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19655_ _19722_/CLK _19655_/D vssd1 vssd1 vccd1 vccd1 _19655_/Q sky130_fd_sc_hd__dfxtp_1
X_16867_ _19347_/Q _16667_/X _16869_/S vssd1 vssd1 vccd1 vccd1 _16868_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18606_ _19553_/CLK _18606_/D vssd1 vssd1 vccd1 vccd1 _18606_/Q sky130_fd_sc_hd__dfxtp_1
X_15818_ _15818_/A vssd1 vssd1 vccd1 vccd1 _18916_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19586_ _19618_/CLK _19586_/D vssd1 vssd1 vccd1 vccd1 _19586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16798_ _16797_/X _19323_/Q _16807_/S vssd1 vssd1 vccd1 vccd1 _16799_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18537_ _18578_/CLK _18537_/D vssd1 vssd1 vccd1 vccd1 _18537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15749_ _15806_/S vssd1 vssd1 vccd1 vccd1 _15758_/S sky130_fd_sc_hd__buf_2
XFILLER_34_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17201__A0 _18444_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09270_ _19078_/Q _11368_/A _11368_/B _11368_/C vssd1 vssd1 vccd1 vccd1 _10857_/B
+ sky130_fd_sc_hd__and4_2
XANTENNA__14015__A0 _18433_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18468_ _19080_/CLK _18468_/D vssd1 vssd1 vccd1 vccd1 _18468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17419_ _17419_/A vssd1 vssd1 vccd1 vccd1 _19576_/D sky130_fd_sc_hd__clkbuf_1
X_18399_ _18401_/CLK _18399_/D vssd1 vssd1 vccd1 vccd1 _18399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12329__A0 _11222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10986__S0 _10668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17245__S _17245_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09552__A _10309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11855__A2 _11820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09606_ _11180_/A _09586_/X _09595_/Y _09605_/Y vssd1 vssd1 vccd1 vccd1 _09606_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_44_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09537_ _10262_/A _09537_/B vssd1 vssd1 vccd1 vccd1 _09537_/X sky130_fd_sc_hd__or2_1
XFILLER_36_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10815__B1 _09177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09468_ _10574_/A _09468_/B vssd1 vssd1 vccd1 vccd1 _09468_/X sky130_fd_sc_hd__or2_1
XFILLER_169_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15754__A0 _14792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_164_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09399_ _10846_/A vssd1 vssd1 vccd1 vccd1 _10589_/A sky130_fd_sc_hd__buf_2
XFILLER_40_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11430_ _11428_/Y _18300_/Q _18299_/Q vssd1 vssd1 vccd1 vccd1 _11430_/X sky130_fd_sc_hd__a21o_1
XFILLER_11_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12137__B _13596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11361_ _11361_/A _11376_/C _13526_/B _13526_/C vssd1 vssd1 vccd1 vccd1 _11366_/A
+ sky130_fd_sc_hd__nor4_4
XFILLER_153_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14633__A _14648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13100_ _18344_/Q _12731_/X _13099_/X _14612_/A vssd1 vssd1 vccd1 vccd1 _18344_/D
+ sky130_fd_sc_hd__o211a_1
X_10312_ _19258_/Q _19029_/Q _18960_/Q _19354_/Q _09701_/S _09555_/X vssd1 vssd1 vccd1
+ vccd1 _10313_/B sky130_fd_sc_hd__mux4_1
XFILLER_98_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14080_ _13949_/A _14079_/X _13950_/X vssd1 vssd1 vccd1 vccd1 _14080_/Y sky130_fd_sc_hd__a21oi_1
X_11292_ _14815_/A vssd1 vssd1 vccd1 vccd1 _14875_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13031_ _13033_/A _13033_/C _13030_/Y vssd1 vssd1 vccd1 vccd1 _18322_/D sky130_fd_sc_hd__o21a_1
X_10243_ _10451_/A _10243_/B vssd1 vssd1 vccd1 vccd1 _10243_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10346__A2 _10335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09831__S1 _09875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input45_A io_ibus_inst[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ _18835_/Q _19389_/Q _19551_/Q _18803_/Q _10131_/S _09610_/X vssd1 vssd1 vccd1
+ vccd1 _10175_/B sky130_fd_sc_hd__mux4_1
XFILLER_160_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14779__S _14893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17770_ _18489_/Q _17770_/B vssd1 vssd1 vccd1 vccd1 _17770_/Y sky130_fd_sc_hd__xnor2_2
X_14982_ _14838_/X _14981_/X _14898_/X vssd1 vssd1 vccd1 vccd1 _14982_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_75_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_89_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16721_ _16721_/A vssd1 vssd1 vccd1 vccd1 _16721_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13933_ _13933_/A vssd1 vssd1 vccd1 vccd1 _14319_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_19440_ _19442_/CLK _19440_/D vssd1 vssd1 vccd1 vccd1 _19440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16652_ _19278_/Q _16651_/X _16655_/S vssd1 vssd1 vccd1 vccd1 _16653_/A sky130_fd_sc_hd__mux2_1
X_13864_ _13864_/A vssd1 vssd1 vccd1 vccd1 _14278_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10401__A _10401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15603_ _18821_/Q _15503_/X _15603_/S vssd1 vssd1 vccd1 vccd1 _15604_/A sky130_fd_sc_hd__mux2_1
X_12815_ _12844_/A _12821_/C vssd1 vssd1 vccd1 vccd1 _12815_/Y sky130_fd_sc_hd__nor2_1
X_19371_ _19534_/CLK _19371_/D vssd1 vssd1 vccd1 vccd1 _19371_/Q sky130_fd_sc_hd__dfxtp_1
X_16583_ _19247_/Q vssd1 vssd1 vccd1 vccd1 _16584_/A sky130_fd_sc_hd__clkbuf_1
X_13795_ _13795_/A vssd1 vssd1 vccd1 vccd1 _13795_/X sky130_fd_sc_hd__clkbuf_2
X_18322_ _19812_/CLK _18322_/D vssd1 vssd1 vccd1 vccd1 _18322_/Q sky130_fd_sc_hd__dfxtp_1
X_15534_ _15534_/A vssd1 vssd1 vccd1 vccd1 _18798_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _18258_/Q vssd1 vssd1 vccd1 vccd1 _12830_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _19855_/CLK _18253_/D vssd1 vssd1 vccd1 vccd1 _18253_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15745__A0 _14753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15465_ _15465_/A vssd1 vssd1 vccd1 vccd1 _18774_/D sky130_fd_sc_hd__clkbuf_1
X_12677_ _18386_/Q _13428_/B _12676_/X vssd1 vssd1 vccd1 vccd1 _12677_/X sky130_fd_sc_hd__a21o_1
XFILLER_129_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17204_ _17204_/A vssd1 vssd1 vccd1 vccd1 _17218_/S sky130_fd_sc_hd__buf_2
XFILLER_31_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14416_ _17751_/A _18516_/Q _14424_/S vssd1 vssd1 vccd1 vccd1 _14417_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18184_ _18249_/A _18184_/B _18185_/B vssd1 vssd1 vccd1 vccd1 _19848_/D sky130_fd_sc_hd__nor3_1
X_11628_ _11628_/A _13524_/C _11628_/C _11517_/X vssd1 vssd1 vccd1 vccd1 _14431_/B
+ sky130_fd_sc_hd__nor4b_4
X_15396_ _15396_/A vssd1 vssd1 vccd1 vccd1 _18745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09975__A1 _09783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17135_ _17135_/A vssd1 vssd1 vccd1 vccd1 _19466_/D sky130_fd_sc_hd__clkbuf_1
X_14347_ _14347_/A vssd1 vssd1 vccd1 vccd1 _18460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11559_ _16212_/D vssd1 vssd1 vccd1 vccd1 _12072_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14543__A _14543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17066_ _17134_/S vssd1 vssd1 vccd1 vccd1 _17075_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_170_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14278_ _14278_/A _14278_/B vssd1 vssd1 vccd1 vccd1 _14278_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14262__B _14265_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16017_ _16017_/A vssd1 vssd1 vccd1 vccd1 _19006_/D sky130_fd_sc_hd__clkbuf_1
X_13229_ _13306_/A vssd1 vssd1 vccd1 vccd1 _13229_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17670__A0 _12727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13287__A1 _19673_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17968_ _19774_/Q _17971_/C _17950_/X vssd1 vssd1 vccd1 vccd1 _17968_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_112_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19707_ _19707_/CLK _19707_/D vssd1 vssd1 vccd1 vccd1 _19707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16919_ _16919_/A _16919_/B _16919_/C vssd1 vssd1 vccd1 vccd1 _17319_/B sky130_fd_sc_hd__and3_1
XFILLER_168_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17899_ _17899_/A vssd1 vssd1 vccd1 vccd1 _19750_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12510__B _12510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19638_ _19638_/CLK _19638_/D vssd1 vssd1 vccd1 vccd1 _19638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19569_ _19569_/CLK _19569_/D vssd1 vssd1 vccd1 vccd1 _19569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16409__S _16413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09889__S1 _09810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09322_ _11056_/A vssd1 vssd1 vccd1 vccd1 _10844_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13622__A _13622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14539__A1 _18564_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09253_ _11497_/A _11519_/A vssd1 vssd1 vccd1 vccd1 _10857_/A sky130_fd_sc_hd__nor2_2
XFILLER_166_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16933__A _16990_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09184_ _09184_/A vssd1 vssd1 vccd1 vccd1 _09712_/A sky130_fd_sc_hd__buf_2
XANTENNA__16144__S _16150_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09718__A1 _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15983__S _15983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09813__S1 _09875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_90_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09577__S0 _09344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17413__A0 _16774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10930_ _10827_/X _10922_/X _10925_/X _10929_/X _09244_/A vssd1 vssd1 vccd1 vccd1
+ _10930_/X sky130_fd_sc_hd__a311o_1
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15975__A0 _14772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10861_ _10548_/X _10860_/X _10871_/A vssd1 vssd1 vccd1 vccd1 _10861_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14628__A _14654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ _12600_/A vssd1 vssd1 vccd1 vccd1 _12600_/X sky130_fd_sc_hd__clkbuf_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13532__A _13532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _13668_/S _13580_/B vssd1 vssd1 vccd1 vccd1 _13712_/B sky130_fd_sc_hd__or2_1
X_10792_ _10634_/X _10788_/X _10790_/X _10899_/A vssd1 vssd1 vccd1 vccd1 _10792_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12531_ _12734_/A _12622_/B vssd1 vssd1 vccd1 vccd1 _12531_/Y sky130_fd_sc_hd__nor2_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12793__D _19856_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ _15250_/A vssd1 vssd1 vccd1 vccd1 _18684_/D sky130_fd_sc_hd__clkbuf_1
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12462_ _12462_/A _12469_/B vssd1 vssd1 vccd1 vccd1 _12462_/Y sky130_fd_sc_hd__nor2_2
XFILLER_138_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14201_ _13978_/X _14203_/B _13979_/X _14200_/X vssd1 vssd1 vccd1 vccd1 _14201_/X
+ sky130_fd_sc_hd__o211a_1
X_11413_ _11413_/A vssd1 vssd1 vccd1 vccd1 _12791_/B sky130_fd_sc_hd__clkbuf_2
X_15181_ _16683_/A vssd1 vssd1 vccd1 vccd1 _15181_/X sky130_fd_sc_hd__buf_2
XFILLER_166_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12393_ _18378_/Q _13388_/A _12393_/C vssd1 vssd1 vccd1 vccd1 _12414_/B sky130_fd_sc_hd__and3_1
XFILLER_4_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14132_ _14054_/X _14122_/X _14131_/Y _14097_/X vssd1 vssd1 vccd1 vccd1 _14132_/X
+ sky130_fd_sc_hd__o211a_1
X_11344_ _11344_/A vssd1 vssd1 vccd1 vccd1 _11375_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09709__A1 _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14063_ _14059_/B _14057_/B _13862_/A _14060_/X _14062_/X vssd1 vssd1 vccd1 vccd1
+ _14063_/X sky130_fd_sc_hd__o221a_1
X_18940_ _19723_/CLK _18940_/D vssd1 vssd1 vccd1 vccd1 _18940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ _11149_/A _11225_/X _11151_/C _11224_/Y _11222_/X vssd1 vssd1 vccd1 vccd1
+ _11275_/Y sky130_fd_sc_hd__o32ai_1
XFILLER_152_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13014_ _13015_/A _13015_/C _18317_/Q vssd1 vssd1 vccd1 vccd1 _13016_/B sky130_fd_sc_hd__a21oi_1
X_10226_ _10226_/A _10226_/B vssd1 vssd1 vccd1 vccd1 _10226_/Y sky130_fd_sc_hd__nor2_1
X_18871_ _19329_/CLK _18871_/D vssd1 vssd1 vccd1 vccd1 _18871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17652__A0 _13245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15194__A _16696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13707__A _13724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17822_ _17822_/A vssd1 vssd1 vccd1 vccd1 _19712_/D sky130_fd_sc_hd__clkbuf_1
X_10157_ _19421_/Q _19197_/Q _19714_/Q _19165_/Q _10154_/S _09146_/A vssd1 vssd1 vccd1
+ vccd1 _10157_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09192__A _19693_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14965_ _14964_/X _18607_/Q _14997_/S vssd1 vssd1 vccd1 vccd1 _14966_/A sky130_fd_sc_hd__mux2_1
X_10088_ _19521_/Q _19135_/Q _19585_/Q _18741_/Q _10114_/S _09769_/A vssd1 vssd1 vccd1
+ vccd1 _10089_/B sky130_fd_sc_hd__mux4_1
X_17753_ _17757_/B _17752_/Y _17713_/X vssd1 vssd1 vccd1 vccd1 _17753_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12330__B _12355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10178__S1 _09610_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16704_ _16704_/A vssd1 vssd1 vccd1 vccd1 _19294_/D sky130_fd_sc_hd__clkbuf_1
X_13916_ _13627_/X _13641_/X _13966_/S vssd1 vssd1 vccd1 vccd1 _13916_/X sky130_fd_sc_hd__mux2_1
X_17684_ _17683_/A _17683_/C _14883_/A vssd1 vssd1 vccd1 vccd1 _17685_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__09893__B1 _09892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14896_ _14969_/A _14912_/B _14896_/C vssd1 vssd1 vccd1 vccd1 _14896_/X sky130_fd_sc_hd__or3_1
XFILLER_62_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19423_ _19810_/CLK _19423_/D vssd1 vssd1 vccd1 vccd1 _19423_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15966__A0 _14729_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16635_ _19273_/Q vssd1 vssd1 vccd1 vccd1 _16636_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__14769__A1 _14768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13847_ _13635_/X _13648_/X _13879_/S vssd1 vssd1 vccd1 vccd1 _13848_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14538__A _16357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16566_ _16566_/A vssd1 vssd1 vccd1 vccd1 _19238_/D sky130_fd_sc_hd__clkbuf_1
X_19354_ _19645_/CLK _19354_/D vssd1 vssd1 vccd1 vccd1 _19354_/Q sky130_fd_sc_hd__dfxtp_1
X_13778_ _13995_/S vssd1 vssd1 vccd1 vccd1 _13838_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18305_ _19790_/CLK _18305_/D vssd1 vssd1 vccd1 vccd1 _18305_/Q sky130_fd_sc_hd__dfxtp_1
X_15517_ _18793_/Q _15516_/X _15520_/S vssd1 vssd1 vccd1 vccd1 _15518_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12729_ _17774_/A _18302_/Q _13090_/S _12728_/X vssd1 vssd1 vccd1 vccd1 _18302_/D
+ sky130_fd_sc_hd__o31a_1
X_19285_ _19285_/CLK _19285_/D vssd1 vssd1 vccd1 vccd1 _19285_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10277__S _10277_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11576__A1_N _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16497_ _16128_/X _19208_/Q _16497_/S vssd1 vssd1 vccd1 vccd1 _16498_/A sky130_fd_sc_hd__mux2_1
X_18236_ _19866_/Q _18232_/B _18235_/Y vssd1 vssd1 vccd1 vccd1 _19866_/D sky130_fd_sc_hd__o21a_1
X_15448_ _18767_/Q _15184_/X _15448_/S vssd1 vssd1 vccd1 vccd1 _15449_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18167_ _19843_/Q _18167_/B vssd1 vssd1 vccd1 vccd1 _18175_/C sky130_fd_sc_hd__and2_1
X_15379_ _15379_/A vssd1 vssd1 vccd1 vccd1 _18737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11755__A1 _19663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17118_ _17118_/A vssd1 vssd1 vccd1 vccd1 _19458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18098_ _18114_/A _18102_/C vssd1 vssd1 vccd1 vccd1 _18098_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12505__B _12505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09940_ _09940_/A _09940_/B _09940_/C vssd1 vssd1 vccd1 vccd1 _09940_/X sky130_fd_sc_hd__or3_4
XFILLER_143_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17049_ _17049_/A vssd1 vssd1 vccd1 vccd1 _17058_/S sky130_fd_sc_hd__buf_4
XFILLER_171_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10306__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09871_ _09942_/A _09871_/B vssd1 vssd1 vccd1 vccd1 _09871_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_112_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14720__B _17391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17643__A0 _19666_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13617__A _13617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14457__A0 _18500_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17523__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15832__A _15878_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11137__A _11137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14209__A0 _18446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11691__A0 _13523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11118__S0 _09583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09305_ _09305_/A vssd1 vssd1 vccd1 vccd1 _09306_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_142_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11443__B1 _11822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09236_ _19660_/Q _19077_/Q _19114_/Q _18720_/Q _09190_/X _09165_/A vssd1 vssd1 vccd1
+ vccd1 _09237_/B sky130_fd_sc_hd__mux4_1
XANTENNA__15185__A1 _15184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13735__A2 _13566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09167_ _10910_/A vssd1 vssd1 vccd1 vccd1 _09168_/A sky130_fd_sc_hd__inv_2
XFILLER_119_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09098_ _11321_/B vssd1 vssd1 vccd1 vccd1 _14519_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11060_ _11060_/A _11060_/B vssd1 vssd1 vccd1 vccd1 _11060_/X sky130_fd_sc_hd__or2_1
XFILLER_88_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12171__A1 _19747_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ _18870_/Q _19328_/Q _10011_/S vssd1 vssd1 vccd1 vccd1 _10011_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09572__C1 _09562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10650__S _10650_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17433__S _17435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14750_ _14765_/C _14745_/Y _14749_/X vssd1 vssd1 vccd1 vccd1 _14750_/Y sky130_fd_sc_hd__o21ai_4
X_11962_ _18361_/Q _18360_/Q _18359_/Q _11962_/D vssd1 vssd1 vccd1 vccd1 _12020_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_44_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13701_ _13761_/A vssd1 vssd1 vccd1 vccd1 _13891_/A sky130_fd_sc_hd__clkbuf_2
X_10913_ _19405_/Q _19181_/Q _19698_/Q _19149_/Q _10909_/X _10910_/X vssd1 vssd1 vccd1
+ vccd1 _10913_/X sky130_fd_sc_hd__mux4_2
XANTENNA__11682__B1 _17241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09970__S0 _09803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14681_ _14578_/A _14633_/X _14680_/X input52/X vssd1 vssd1 vccd1 vccd1 _14682_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16049__S _16049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11893_ _11940_/A vssd1 vssd1 vccd1 vccd1 _12057_/A sky130_fd_sc_hd__buf_2
X_16420_ _19174_/Q _15577_/X _16424_/S vssd1 vssd1 vccd1 vccd1 _16421_/A sky130_fd_sc_hd__mux2_1
X_13632_ _13682_/S vssd1 vssd1 vccd1 vccd1 _13659_/S sky130_fd_sc_hd__clkbuf_2
X_10844_ _10844_/A _10844_/B vssd1 vssd1 vccd1 vccd1 _10844_/X sky130_fd_sc_hd__or2_1
XANTENNA__09627__B1 _09625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13423__B2 _18649_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16351_ _16128_/X _19144_/Q _16351_/S vssd1 vssd1 vccd1 vccd1 _16352_/A sky130_fd_sc_hd__mux2_1
X_13563_ _13563_/A _13563_/B vssd1 vssd1 vccd1 vccd1 _13564_/A sky130_fd_sc_hd__and2_1
XFILLER_158_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10775_ _10769_/Y _10771_/X _10773_/X _10946_/A _10774_/X vssd1 vssd1 vccd1 vccd1
+ _10780_/B sky130_fd_sc_hd__o221a_1
XFILLER_40_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10332__S1 _09735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15302_ _15324_/A vssd1 vssd1 vccd1 vccd1 _15311_/S sky130_fd_sc_hd__clkbuf_4
X_19070_ _19718_/CLK _19070_/D vssd1 vssd1 vccd1 vccd1 _19070_/Q sky130_fd_sc_hd__dfxtp_1
X_12514_ _13171_/A _18635_/Q vssd1 vssd1 vccd1 vccd1 _12514_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16282_ _16282_/A vssd1 vssd1 vccd1 vccd1 _19113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13494_ _13494_/A vssd1 vssd1 vccd1 vccd1 _18405_/D sky130_fd_sc_hd__clkbuf_1
X_18021_ _18023_/A _18023_/B _17993_/X vssd1 vssd1 vccd1 vccd1 _18021_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_74_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15233_ _18680_/Q _15232_/X _15233_/S vssd1 vssd1 vccd1 vccd1 _15234_/A sky130_fd_sc_hd__mux2_1
X_12445_ _14332_/B _12446_/B vssd1 vssd1 vccd1 vccd1 _14331_/A sky130_fd_sc_hd__nand2_1
XFILLER_173_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14093__A _14093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11737__A1 _18565_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11510__A _13523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09187__A _10107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15164_ _15164_/A vssd1 vssd1 vccd1 vccd1 _18658_/D sky130_fd_sc_hd__clkbuf_1
X_12376_ _11517_/B _13525_/A _12345_/X _12502_/A vssd1 vssd1 vccd1 vccd1 _12377_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14115_ _14115_/A vssd1 vssd1 vccd1 vccd1 _14115_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11327_ _18582_/Q vssd1 vssd1 vccd1 vccd1 _11514_/A sky130_fd_sc_hd__buf_2
XANTENNA__16512__S _16514_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15095_ _15095_/A _15095_/B vssd1 vssd1 vccd1 vccd1 _15125_/A sky130_fd_sc_hd__nor2_2
XFILLER_107_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09789__S0 _09760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18923_ _19707_/CLK _18923_/D vssd1 vssd1 vccd1 vccd1 _18923_/Q sky130_fd_sc_hd__dfxtp_1
X_14046_ _13942_/A _14043_/Y _14045_/Y _13711_/B vssd1 vssd1 vccd1 vccd1 _14046_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA_output76_A _11978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11258_ _11258_/A _11258_/B _11258_/C _10979_/X vssd1 vssd1 vccd1 vccd1 _11258_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17625__A0 _19663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09563__C1 _09562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13437__A _15262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10209_ _19646_/Q _19063_/Q _19100_/Q _18706_/Q _09795_/A _10080_/X vssd1 vssd1 vccd1
+ vccd1 _10210_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12341__A _18376_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18854_ _19569_/CLK _18854_/D vssd1 vssd1 vccd1 vccd1 _18854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14032__S _14032_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11189_ _11189_/A _11189_/B vssd1 vssd1 vccd1 vccd1 _11189_/Y sky130_fd_sc_hd__nand2_1
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17805_ _15168_/X _19705_/Q _17805_/S vssd1 vssd1 vccd1 vccd1 _17806_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15100__A1 _18626_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18785_ _19534_/CLK _18785_/D vssd1 vssd1 vccd1 vccd1 _18785_/Q sky130_fd_sc_hd__dfxtp_1
X_15997_ _14889_/X _18997_/Q _16005_/S vssd1 vssd1 vccd1 vccd1 _15998_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17736_ _17736_/A vssd1 vssd1 vccd1 vccd1 _19682_/D sky130_fd_sc_hd__clkbuf_1
X_14948_ input13/X _14924_/X _14925_/X vssd1 vssd1 vccd1 vccd1 _14948_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09961__S0 _09803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14879_ _16790_/A vssd1 vssd1 vccd1 vccd1 _14879_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17667_ _18469_/Q _18470_/Q _17667_/C vssd1 vssd1 vccd1 vccd1 _17674_/B sky130_fd_sc_hd__or3_1
XFILLER_165_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19406_ _19699_/CLK _19406_/D vssd1 vssd1 vccd1 vccd1 _19406_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10571__S1 _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16618_ _16618_/A vssd1 vssd1 vccd1 vccd1 _19264_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17598_ _17598_/A vssd1 vssd1 vccd1 vccd1 _19656_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15798__S _15802_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16549_ _16560_/A vssd1 vssd1 vccd1 vccd1 _16558_/S sky130_fd_sc_hd__buf_4
XANTENNA__09713__S0 _10257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19337_ _19337_/CLK _19337_/D vssd1 vssd1 vccd1 vccd1 _19337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19268_ _19331_/CLK _19268_/D vssd1 vssd1 vccd1 vccd1 _19268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18219_ _19861_/Q _18222_/C vssd1 vssd1 vccd1 vccd1 _18221_/A sky130_fd_sc_hd__and2_1
XFILLER_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19199_ _19810_/CLK _19199_/D vssd1 vssd1 vccd1 vccd1 _19199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12516__A _12516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17518__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17864__B1 _14638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16422__S _16424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09923_ _09278_/X _09910_/X _09922_/X _09285_/X _18449_/Q vssd1 vssd1 vccd1 vccd1
+ _09951_/A sky130_fd_sc_hd__a32o_4
XANTENNA__12153__A1 _11997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09854_ _09854_/A _09854_/B _09854_/C vssd1 vssd1 vccd1 vccd1 _09854_/X sky130_fd_sc_hd__or3_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11900__A1 _11901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10703__A2 _10702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _09905_/A _09784_/X _09231_/A vssd1 vssd1 vccd1 vccd1 _09785_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16658__A _16741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14850__A0 _18438_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13405__B2 _18379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11967__A1 _14543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10560_ _18858_/Q _19316_/Q _10560_/S vssd1 vssd1 vccd1 vccd1 _10560_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13169__B1 _14673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ _19434_/Q _19210_/Q _19727_/Q _19178_/Q _09190_/X _09165_/A vssd1 vssd1 vccd1
+ vccd1 _09219_/X sky130_fd_sc_hd__mux4_2
XANTENNA__14905__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10491_ _18764_/Q _18993_/Q _18924_/Q _19222_/Q _09522_/A _10238_/A vssd1 vssd1 vccd1
+ vccd1 _10492_/B sky130_fd_sc_hd__mux4_1
X_12230_ _14227_/A _12230_/B vssd1 vssd1 vccd1 vccd1 _12233_/A sky130_fd_sc_hd__xnor2_2
XFILLER_136_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12392__A1 _13388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12161_ _12161_/A _12161_/B vssd1 vssd1 vccd1 vccd1 _12163_/A sky130_fd_sc_hd__nor2_2
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16332__S _16340_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11112_ _18599_/Q _19288_/Q _11112_/S vssd1 vssd1 vccd1 vccd1 _11113_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11984__B _19739_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09735__A _09735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12092_ _12095_/A _12092_/B vssd1 vssd1 vccd1 vccd1 _12092_/X sky130_fd_sc_hd__or2_1
XFILLER_2_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11043_ _10996_/A _11042_/X _09223_/A vssd1 vssd1 vccd1 vccd1 _11043_/Y sky130_fd_sc_hd__o21ai_1
X_15920_ _14918_/X _18962_/Q _15924_/S vssd1 vssd1 vccd1 vccd1 _15921_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10155__B1 _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15851_ _15851_/A vssd1 vssd1 vccd1 vccd1 _18931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14802_ _14802_/A _14802_/B _14900_/A input30/X vssd1 vssd1 vccd1 vccd1 _14803_/B
+ sky130_fd_sc_hd__and4_1
X_15782_ _15793_/A vssd1 vssd1 vccd1 vccd1 _15791_/S sky130_fd_sc_hd__buf_4
X_18570_ _18578_/CLK _18570_/D vssd1 vssd1 vccd1 vccd1 _18570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12994_ _13034_/A _12994_/B _12994_/C vssd1 vssd1 vccd1 vccd1 _18311_/D sky130_fd_sc_hd__nor3_1
XANTENNA__13644__A1 _12446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11104__C1 _09246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10458__A1 _09402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17521_ _19622_/Q _16721_/X _17529_/S vssd1 vssd1 vccd1 vccd1 _17522_/A sky130_fd_sc_hd__mux2_1
X_14733_ _19081_/Q vssd1 vssd1 vccd1 vccd1 _14873_/A sky130_fd_sc_hd__inv_2
XANTENNA__09943__S0 _09866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11945_ _12478_/B _11831_/X _12023_/B _11944_/Y vssd1 vssd1 vccd1 vccd1 _12030_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _17452_/A vssd1 vssd1 vccd1 vccd1 _19591_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _14672_/A _15952_/B vssd1 vssd1 vccd1 vccd1 _18574_/D sky130_fd_sc_hd__nor2_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _11842_/A _13658_/A _11875_/X vssd1 vssd1 vccd1 vccd1 _11876_/X sky130_fd_sc_hd__o21a_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16403_ _16403_/A vssd1 vssd1 vccd1 vccd1 _19166_/D sky130_fd_sc_hd__clkbuf_1
X_13615_ _13615_/A vssd1 vssd1 vccd1 vccd1 _13615_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17383_ _16835_/X _19561_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _17384_/A sky130_fd_sc_hd__mux2_1
X_10827_ _10827_/A vssd1 vssd1 vccd1 vccd1 _10827_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14595_ _11297_/C _12731_/A _14593_/X _14594_/Y vssd1 vssd1 vccd1 vccd1 _14596_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16334_ _16103_/X _19136_/Q _16340_/S vssd1 vssd1 vccd1 vccd1 _16335_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13720__A _13720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19122_ _19614_/CLK _19122_/D vssd1 vssd1 vccd1 vccd1 _19122_/Q sky130_fd_sc_hd__dfxtp_1
X_13546_ _13521_/X _13522_/X _13545_/X _14516_/S vssd1 vssd1 vccd1 vccd1 _13546_/X
+ sky130_fd_sc_hd__a31o_1
X_10758_ _09274_/A _10748_/X _10757_/X _09281_/A _18432_/Q vssd1 vssd1 vccd1 vccd1
+ _11075_/A sky130_fd_sc_hd__a32o_2
XFILLER_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19053_ _19614_/CLK _19053_/D vssd1 vssd1 vccd1 vccd1 _19053_/Q sky130_fd_sc_hd__dfxtp_1
X_16265_ _16265_/A vssd1 vssd1 vccd1 vccd1 _19105_/D sky130_fd_sc_hd__clkbuf_1
X_13477_ _13499_/A vssd1 vssd1 vccd1 vccd1 _13486_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__10630__B2 _18434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10689_ _09179_/A _10688_/X _09224_/A vssd1 vssd1 vccd1 vccd1 _10689_/X sky130_fd_sc_hd__o21a_1
X_15216_ _16718_/A vssd1 vssd1 vccd1 vccd1 _15216_/X sky130_fd_sc_hd__clkbuf_2
X_18004_ _19786_/Q _18006_/C _18003_/Y vssd1 vssd1 vccd1 vccd1 _19786_/D sky130_fd_sc_hd__o21a_1
XANTENNA__10069__S0 _10033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12428_ _12428_/A vssd1 vssd1 vccd1 vccd1 _12430_/A sky130_fd_sc_hd__inv_2
XFILLER_138_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16196_ _16196_/A vssd1 vssd1 vccd1 vccd1 _16205_/S sky130_fd_sc_hd__buf_6
XFILLER_126_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15147_ _18653_/Q _15146_/X _15153_/S vssd1 vssd1 vccd1 vccd1 _15148_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12359_ _19755_/Q vssd1 vssd1 vccd1 vccd1 _12361_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__16242__S _16246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15078_ _15078_/A vssd1 vssd1 vccd1 vccd1 _18617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13167__A _17781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18906_ _19554_/CLK _18906_/D vssd1 vssd1 vccd1 vccd1 _18906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14029_ _14314_/A _14020_/X _14028_/X _14054_/A vssd1 vssd1 vccd1 vccd1 _14029_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12071__A _19674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10146__B1 _09621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18837_ _19553_/CLK _18837_/D vssd1 vssd1 vccd1 vccd1 _18837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17073__S _17075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09570_ _19626_/Q _19464_/Q _18910_/Q _18680_/Q _09700_/A _09642_/A vssd1 vssd1 vccd1
+ vccd1 _09571_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09839__B1 _09625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18768_ _19551_/CLK _18768_/D vssd1 vssd1 vccd1 vccd1 _18768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09934__S0 _09866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17719_ _17719_/A vssd1 vssd1 vccd1 vccd1 _19679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18699_ _19706_/CLK _18699_/D vssd1 vssd1 vccd1 vccd1 _18699_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17801__S _17805_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13333__C _14958_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13630__A _13630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10465__S _10465_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12246__A _12246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14902__A4 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_clock_A clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09555__A _09642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09906_ _19620_/Q _19458_/Q _18904_/Q _18674_/Q _09782_/X _09783_/X vssd1 vssd1 vccd1
+ vccd1 _09906_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13874__A1 _11667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09837_ _09320_/X _09819_/Y _09830_/X _09836_/Y _09395_/X vssd1 vssd1 vccd1 vccd1
+ _09837_/X sky130_fd_sc_hd__o311a_4
XFILLER_100_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10232__S0 _10230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09768_ _10103_/A vssd1 vssd1 vccd1 vccd1 _09769_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09699_ _18612_/Q _19301_/Q _10256_/S vssd1 vssd1 vccd1 vccd1 _09699_/X sky130_fd_sc_hd__mux2_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11325__A _14578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11730_ _15262_/A _11728_/X _11801_/A vssd1 vssd1 vccd1 vccd1 _11730_/X sky130_fd_sc_hd__a21o_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _17221_/A vssd1 vssd1 vccd1 vccd1 _17143_/S sky130_fd_sc_hd__clkbuf_4
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16327__S _16329_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13400_ _18378_/Q _13413_/B vssd1 vssd1 vccd1 vccd1 _13400_/X sky130_fd_sc_hd__or2_1
X_10612_ _19693_/Q vssd1 vssd1 vccd1 vccd1 _10992_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_168_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14380_ _18472_/Q vssd1 vssd1 vccd1 vccd1 _17683_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11592_ _11592_/A vssd1 vssd1 vccd1 vccd1 _12259_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_128_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13331_ _18324_/Q _13178_/X _12749_/X _19813_/Q vssd1 vssd1 vccd1 vccd1 _13331_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10543_ _09442_/X _10540_/X _10542_/X vssd1 vssd1 vccd1 vccd1 _10543_/X sky130_fd_sc_hd__a21o_1
X_16050_ _16050_/A vssd1 vssd1 vccd1 vccd1 _19018_/D sky130_fd_sc_hd__clkbuf_1
X_13262_ _13185_/X _13259_/X _13261_/X _13232_/X vssd1 vssd1 vccd1 vccd1 _18360_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10474_ _19640_/Q _19057_/Q _19094_/Q _18700_/Q _09631_/A _09635_/A vssd1 vssd1 vccd1
+ vccd1 _10475_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12365__A1 _19686_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_160_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19534_/CLK sky130_fd_sc_hd__clkbuf_16
X_15001_ input18/X _14960_/X _15000_/X vssd1 vssd1 vccd1 vccd1 _15001_/X sky130_fd_sc_hd__a21o_1
XFILLER_124_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12213_ _14211_/A vssd1 vssd1 vccd1 vccd1 _12213_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13193_ _19861_/Q _12604_/A _12583_/A _18131_/B vssd1 vssd1 vccd1 vccd1 _13193_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16062__S _16065_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12144_ _19745_/Q _19746_/Q _12144_/C vssd1 vssd1 vccd1 vccd1 _12215_/C sky130_fd_sc_hd__and3_1
XANTENNA__09465__A _11097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15303__A1 _15187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_clock_A clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16997__S _17003_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19740_ _19753_/CLK _19740_/D vssd1 vssd1 vccd1 vccd1 _19740_/Q sky130_fd_sc_hd__dfxtp_1
X_12075_ _18365_/Q _18364_/Q _12075_/C vssd1 vssd1 vccd1 vccd1 _12123_/C sky130_fd_sc_hd__and3_2
XFILLER_111_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16952_ _16952_/A vssd1 vssd1 vccd1 vccd1 _19384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_175_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19704_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_6_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_159_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11026_ _11026_/A _11026_/B vssd1 vssd1 vccd1 vccd1 _11026_/Y sky130_fd_sc_hd__nor2_1
X_15903_ _15903_/A vssd1 vssd1 vccd1 vccd1 _18954_/D sky130_fd_sc_hd__clkbuf_1
X_19671_ _19687_/CLK _19671_/D vssd1 vssd1 vccd1 vccd1 _19671_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_65_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16883_ _19354_/Q _16689_/X _16891_/S vssd1 vssd1 vccd1 vccd1 _16884_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16298__A _16355_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13715__A _14274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18622_ _19468_/CLK _18622_/D vssd1 vssd1 vccd1 vccd1 _18622_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__15406__S _15406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15834_ _15834_/A vssd1 vssd1 vccd1 vccd1 _18923_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14814__B1 _14813_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18553_ _18564_/CLK _18553_/D vssd1 vssd1 vccd1 vccd1 _18553_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ _18306_/Q _12973_/C _12976_/Y vssd1 vssd1 vccd1 vccd1 _18306_/D sky130_fd_sc_hd__o21a_1
X_15765_ _14856_/X _18893_/Q _15769_/S vssd1 vssd1 vccd1 vccd1 _15766_/A sky130_fd_sc_hd__mux2_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17504_ _17504_/A vssd1 vssd1 vccd1 vccd1 _19614_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11928_ _12152_/B vssd1 vssd1 vccd1 vccd1 _11928_/X sky130_fd_sc_hd__clkbuf_2
X_14716_ _14716_/A vssd1 vssd1 vccd1 vccd1 _16919_/B sky130_fd_sc_hd__clkbuf_1
X_18484_ _18487_/CLK _18484_/D vssd1 vssd1 vccd1 vccd1 _18484_/Q sky130_fd_sc_hd__dfxtp_1
X_15696_ _15696_/A vssd1 vssd1 vccd1 vccd1 _18862_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17435_ _16806_/X _19584_/Q _17435_/S vssd1 vssd1 vccd1 vccd1 _17436_/A sky130_fd_sc_hd__mux2_1
X_14647_ _14672_/A _17774_/B vssd1 vssd1 vccd1 vccd1 _18569_/D sky130_fd_sc_hd__nor2_1
XFILLER_162_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11859_ _12152_/B vssd1 vssd1 vccd1 vccd1 _11859_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14042__A1 _14126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_113_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19738_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_82_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15141__S _15153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13250__C1 _13249_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17366_ _16809_/X _19553_/Q _17374_/S vssd1 vssd1 vccd1 vccd1 _17367_/A sky130_fd_sc_hd__mux2_1
X_14578_ _14578_/A _14580_/B vssd1 vssd1 vccd1 vccd1 _14578_/X sky130_fd_sc_hd__or2_1
XFILLER_174_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14265__B _14265_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19105_ _19718_/CLK _19105_/D vssd1 vssd1 vccd1 vccd1 _19105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17857__A _17890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16317_ _16317_/A vssd1 vssd1 vccd1 vccd1 _19128_/D sky130_fd_sc_hd__clkbuf_1
X_13529_ _13529_/A _13529_/B _13587_/A _13529_/D vssd1 vssd1 vccd1 vccd1 _13529_/X
+ sky130_fd_sc_hd__and4_1
X_17297_ _17297_/A vssd1 vssd1 vccd1 vccd1 _19522_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19036_ _19838_/CLK _19036_/D vssd1 vssd1 vccd1 vccd1 _19036_/Q sky130_fd_sc_hd__dfxtp_1
X_16248_ _16270_/A vssd1 vssd1 vccd1 vccd1 _16257_/S sky130_fd_sc_hd__buf_2
XFILLER_134_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_128_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _18482_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_173_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17819__A0 _15187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput103 _11880_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[8] sky130_fd_sc_hd__buf_2
Xoutput114 _12480_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[12] sky130_fd_sc_hd__buf_2
X_16179_ _16090_/X _19063_/Q _16183_/S vssd1 vssd1 vccd1 vccd1 _16180_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput125 _12494_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[22] sky130_fd_sc_hd__buf_2
Xoutput136 _12464_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[3] sky130_fd_sc_hd__buf_2
Xoutput147 _12003_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[12] sky130_fd_sc_hd__buf_2
XFILLER_99_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput158 _17898_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[22] sky130_fd_sc_hd__buf_2
XFILLER_82_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput169 _17860_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[3] sky130_fd_sc_hd__buf_2
XFILLER_141_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17592__A _17592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16700__S _16703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10214__S0 _09545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11129__B _12481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19869_ _19871_/CLK _19869_/D vssd1 vssd1 vccd1 vccd1 _19869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15316__S _15322_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10765__S1 _09482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09622_ _10182_/A _09620_/X _09621_/X vssd1 vssd1 vccd1 vccd1 _09622_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_28_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09907__S0 _09976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _09643_/S vssd1 vssd1 vccd1 vccd1 _09553_/X sky130_fd_sc_hd__buf_4
XANTENNA__14281__A1 _12333_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17531__S _17533_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11095__A1 _09434_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09484_ _19273_/Q _19044_/Q _18975_/Q _19369_/Q _10389_/S _09483_/X vssd1 vssd1 vccd1
+ vccd1 _09485_/B sky130_fd_sc_hd__mux4_1
XFILLER_51_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_92_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19855_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_133_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10453__S0 _10224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10190_ _11178_/A _10189_/X _09317_/A vssd1 vssd1 vccd1 vccd1 _10190_/X sky130_fd_sc_hd__o21a_1
XFILLER_87_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_160_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10205__S0 _09545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12900_ _12910_/D _12897_/B _12869_/X vssd1 vssd1 vccd1 vccd1 _12900_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_46_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13880_ _13757_/X _13765_/X _13880_/S vssd1 vssd1 vccd1 vccd1 _13993_/B sky130_fd_sc_hd__mux2_1
XFILLER_100_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12831_ _12851_/A _12831_/B _12831_/C vssd1 vssd1 vccd1 vccd1 _18259_/D sky130_fd_sc_hd__nor3_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _15550_/A vssd1 vssd1 vccd1 vccd1 _18803_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_30_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19584_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _14565_/A vssd1 vssd1 vccd1 vccd1 _14519_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14501_/A vssd1 vssd1 vccd1 vccd1 _18520_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11713_ _11706_/X _11709_/X _11711_/X _12696_/A vssd1 vssd1 vccd1 vccd1 _11713_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15481_ _18782_/Q _15232_/X _15481_/S vssd1 vssd1 vccd1 vccd1 _15482_/A sky130_fd_sc_hd__mux2_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _13104_/B _12661_/X _12689_/X _12692_/X vssd1 vssd1 vccd1 vccd1 _18335_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _17220_/A vssd1 vssd1 vccd1 vccd1 _19492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _19468_/D _14432_/B vssd1 vssd1 vccd1 vccd1 _14591_/B sky130_fd_sc_hd__nor2_4
X_11644_ _11644_/A _11644_/B vssd1 vssd1 vccd1 vccd1 _13571_/C sky130_fd_sc_hd__nor2_1
XFILLER_168_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17151_ _19472_/Q _17150_/X _17155_/S vssd1 vssd1 vccd1 vccd1 _17152_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15896__S _15902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19622_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14363_ _18466_/Q vssd1 vssd1 vccd1 vccd1 _17645_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_85_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11575_ _11692_/A _11575_/B _15095_/B vssd1 vssd1 vccd1 vccd1 _11575_/Y sky130_fd_sc_hd__nor3_1
Xinput16 io_dbus_rdata[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_2
Xinput27 io_dbus_rdata[4] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_2
X_16102_ _16102_/A vssd1 vssd1 vccd1 vccd1 _19034_/D sky130_fd_sc_hd__clkbuf_1
X_13314_ _18367_/Q _13319_/B vssd1 vssd1 vccd1 vccd1 _13314_/X sky130_fd_sc_hd__or2_1
Xinput38 io_ibus_inst[13] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_2
Xinput49 io_ibus_inst[23] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_2
X_17082_ _16768_/X _19442_/Q _17086_/S vssd1 vssd1 vccd1 vccd1 _17083_/A sky130_fd_sc_hd__mux2_1
X_10526_ _09679_/A _10525_/X _09314_/A vssd1 vssd1 vccd1 vccd1 _10526_/X sky130_fd_sc_hd__o21a_1
XFILLER_128_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14294_ _13909_/X _14292_/X _14293_/Y _15123_/A vssd1 vssd1 vccd1 vccd1 _14294_/X
+ sky130_fd_sc_hd__a31o_1
X_16033_ _16743_/A vssd1 vssd1 vccd1 vccd1 _16033_/X sky130_fd_sc_hd__clkbuf_1
X_13245_ _13217_/X _13234_/Y _13244_/X _13229_/X _18628_/Q vssd1 vssd1 vccd1 vccd1
+ _13245_/X sky130_fd_sc_hd__a32o_4
XANTENNA__15197__A _16699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10457_ _09681_/X _10447_/Y _10452_/X _10456_/Y _09393_/A vssd1 vssd1 vccd1 vccd1
+ _10457_/X sky130_fd_sc_hd__o311a_1
XFILLER_6_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09195__A _10875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ _19796_/Q vssd1 vssd1 vccd1 vccd1 _18031_/B sky130_fd_sc_hd__clkbuf_2
X_10388_ _10388_/A vssd1 vssd1 vccd1 vccd1 _10388_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10995__S1 _10960_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ _14557_/A _12026_/X _12226_/A _12487_/A vssd1 vssd1 vccd1 vccd1 _12128_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_151_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17984_ _19780_/Q _17988_/C _17950_/X vssd1 vssd1 vccd1 vccd1 _17984_/Y sky130_fd_sc_hd__a21oi_1
X_19723_ _19723_/CLK _19723_/D vssd1 vssd1 vccd1 vccd1 _19723_/Q sky130_fd_sc_hd__dfxtp_1
X_16935_ _16935_/A vssd1 vssd1 vccd1 vccd1 _19376_/D sky130_fd_sc_hd__clkbuf_1
X_12058_ _12131_/A _12131_/B _12348_/A vssd1 vssd1 vccd1 vccd1 _12059_/B sky130_fd_sc_hd__o21ai_1
XFILLER_77_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11009_ _18754_/Q _18983_/Q _18914_/Q _19212_/Q _18977_/Q _18978_/Q vssd1 vssd1 vccd1
+ vccd1 _11010_/B sky130_fd_sc_hd__mux4_1
XFILLER_42_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19654_ _19657_/CLK _19654_/D vssd1 vssd1 vccd1 vccd1 _19654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_6_0_clock_A clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16866_ _16866_/A vssd1 vssd1 vccd1 vccd1 _19346_/D sky130_fd_sc_hd__clkbuf_1
X_18605_ _19716_/CLK _18605_/D vssd1 vssd1 vccd1 vccd1 _18605_/Q sky130_fd_sc_hd__dfxtp_1
X_15817_ _14753_/X _18916_/Q _15819_/S vssd1 vssd1 vccd1 vccd1 _15818_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19585_ _19716_/CLK _19585_/D vssd1 vssd1 vccd1 vccd1 _19585_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14263__A1 _11602_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16797_ _16797_/A vssd1 vssd1 vccd1 vccd1 _16797_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12274__B1 _17693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18536_ _18567_/CLK _18536_/D vssd1 vssd1 vccd1 vccd1 _18536_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ _15748_/A vssd1 vssd1 vccd1 vccd1 _18885_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17201__A1 _12617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18467_ _18632_/CLK _18467_/D vssd1 vssd1 vccd1 vccd1 _18467_/Q sky130_fd_sc_hd__dfxtp_1
X_15679_ _15679_/A vssd1 vssd1 vccd1 vccd1 _18854_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17418_ _16781_/X _19576_/Q _17424_/S vssd1 vssd1 vccd1 vccd1 _17419_/A sky130_fd_sc_hd__mux2_1
X_18398_ _19690_/CLK _18398_/D vssd1 vssd1 vccd1 vccd1 _18398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17349_ _17349_/A vssd1 vssd1 vccd1 vccd1 _19545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11805__A1_N _12468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10309__A _10309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14318__A2 _13873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12329__A1 _18516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19019_ _19634_/CLK _19019_/D vssd1 vssd1 vccd1 vccd1 _19019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12524__A _12603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10986__S1 _10906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13829__A1 _11624_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18211__A _18214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10512__B1 _10593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09605_ _10325_/A _09604_/X _09616_/A vssd1 vssd1 vccd1 vccd1 _09605_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_16_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17261__S _17269_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09536_ _19272_/Q _19043_/Q _18974_/Q _19368_/Q _11157_/S _09144_/A vssd1 vssd1 vccd1
+ vccd1 _09537_/B sky130_fd_sc_hd__mux4_1
XFILLER_25_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11068__B2 _11046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10815__A1 _09169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09467_ _19627_/Q _19465_/Q _18911_/Q _18681_/Q _10540_/S _09141_/A vssd1 vssd1 vccd1
+ vccd1 _09468_/B sky130_fd_sc_hd__mux4_1
XFILLER_24_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_107_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09398_ _10944_/A vssd1 vssd1 vccd1 vccd1 _10846_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11360_ _11477_/A _11587_/A _11360_/C _11587_/B vssd1 vssd1 vccd1 vccd1 _11367_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10311_ _09214_/A _10302_/X _10305_/X _10310_/X _09247_/A vssd1 vssd1 vccd1 vccd1
+ _10311_/X sky130_fd_sc_hd__a311o_2
XFILLER_164_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11291_ _19079_/Q vssd1 vssd1 vccd1 vccd1 _14815_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12434__A _19758_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13030_ _13033_/A _13033_/C _13011_/X vssd1 vssd1 vccd1 vccd1 _13030_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10242_ _18603_/Q _19292_/Q _10242_/S vssd1 vssd1 vccd1 vccd1 _10243_/B sky130_fd_sc_hd__mux2_1
XFILLER_133_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09951__B_N _12495_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10346__A3 _10344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16340__S _16340_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10173_ _10182_/A _10173_/B vssd1 vssd1 vccd1 vccd1 _10173_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18121__A _18199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input38_A io_ibus_inst[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14981_ _18449_/Q _12756_/B _14981_/S vssd1 vssd1 vccd1 vccd1 _14981_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13296__A2 _13294_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_opt_5_0_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_5_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
X_16720_ _16720_/A vssd1 vssd1 vccd1 vccd1 _19299_/D sky130_fd_sc_hd__clkbuf_1
X_13932_ _13738_/X _13918_/X _13931_/X _13909_/X vssd1 vssd1 vccd1 vccd1 _13932_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16651_ _16651_/A vssd1 vssd1 vccd1 vccd1 _16651_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13863_ _13863_/A vssd1 vssd1 vccd1 vccd1 _13864_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12814_ _12823_/D vssd1 vssd1 vccd1 vccd1 _12821_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15602_ _15602_/A vssd1 vssd1 vccd1 vccd1 _18820_/D sky130_fd_sc_hd__clkbuf_1
X_19370_ _19628_/CLK _19370_/D vssd1 vssd1 vccd1 vccd1 _19370_/Q sky130_fd_sc_hd__dfxtp_1
X_16582_ _16582_/A vssd1 vssd1 vccd1 vccd1 _19246_/D sky130_fd_sc_hd__clkbuf_1
X_13794_ _13856_/A vssd1 vssd1 vccd1 vccd1 _13795_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18321_ _19810_/CLK _18321_/D vssd1 vssd1 vccd1 vccd1 _18321_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11154__S1 _10306_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12745_ _19682_/Q _12737_/X _12740_/X _12744_/X vssd1 vssd1 vccd1 vccd1 _12745_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__17195__A0 _18442_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15533_ _18798_/Q _15532_/X _15536_/S vssd1 vssd1 vccd1 vccd1 _15534_/A sky130_fd_sc_hd__mux2_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11513__A _11513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18252_ _19872_/CLK _18252_/D vssd1 vssd1 vccd1 vccd1 _18252_/Q sky130_fd_sc_hd__dfxtp_1
X_15464_ _18774_/Q _15207_/X _15470_/S vssd1 vssd1 vccd1 vccd1 _15465_/A sky130_fd_sc_hd__mux2_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _18335_/Q _12564_/A _12606_/A _12873_/B _12641_/A vssd1 vssd1 vccd1 vccd1
+ _12676_/X sky130_fd_sc_hd__a221o_1
XANTENNA__16942__A0 _16774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17203_ _17203_/A vssd1 vssd1 vccd1 vccd1 _19487_/D sky130_fd_sc_hd__clkbuf_1
X_14415_ _18484_/Q vssd1 vssd1 vccd1 vccd1 _17751_/A sky130_fd_sc_hd__clkbuf_2
X_11627_ _17611_/B vssd1 vssd1 vccd1 vccd1 _12715_/B sky130_fd_sc_hd__clkbuf_4
X_18183_ _19848_/Q _19847_/Q _18183_/C vssd1 vssd1 vccd1 vccd1 _18185_/B sky130_fd_sc_hd__and3_1
X_15395_ _18745_/Q _15216_/X _15395_/S vssd1 vssd1 vccd1 vccd1 _15396_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09424__A1 _09415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17134_ _16844_/X _19466_/Q _17134_/S vssd1 vssd1 vccd1 vccd1 _17135_/A sky130_fd_sc_hd__mux2_1
X_14346_ _14743_/A _18492_/Q _14352_/S vssd1 vssd1 vccd1 vccd1 _14347_/A sky130_fd_sc_hd__mux2_1
X_11558_ _14718_/B vssd1 vssd1 vccd1 vccd1 _16212_/D sky130_fd_sc_hd__buf_4
XFILLER_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17065_ _17121_/A vssd1 vssd1 vccd1 vccd1 _17134_/S sky130_fd_sc_hd__buf_6
X_10509_ _18859_/Q _19317_/Q _10581_/S vssd1 vssd1 vccd1 vccd1 _10510_/B sky130_fd_sc_hd__mux2_1
X_14277_ _14274_/B _14272_/B _13856_/A _14275_/X _14276_/X vssd1 vssd1 vccd1 vccd1
+ _14278_/B sky130_fd_sc_hd__o221a_1
X_11489_ _11282_/A _11585_/A _11485_/A _14547_/A vssd1 vssd1 vccd1 vccd1 _15079_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16016_ _14996_/X _19006_/Q _16016_/S vssd1 vssd1 vccd1 vccd1 _16017_/A sky130_fd_sc_hd__mux2_1
X_13228_ _18627_/Q _13228_/B vssd1 vssd1 vccd1 vccd1 _13228_/X sky130_fd_sc_hd__or2_1
XANTENNA__10933__A_N _09481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12063__B _13603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17346__S _17352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _19762_/Q vssd1 vssd1 vccd1 vccd1 _17934_/B sky130_fd_sc_hd__clkbuf_2
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _19773_/Q _17965_/B _17966_/Y vssd1 vssd1 vccd1 vccd1 _19773_/D sky130_fd_sc_hd__o21a_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13287__A2 _12668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19706_ _19706_/CLK _19706_/D vssd1 vssd1 vccd1 vccd1 _19706_/Q sky130_fd_sc_hd__dfxtp_1
X_16918_ _16918_/A vssd1 vssd1 vccd1 vccd1 _19370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17898_ _17909_/A _17898_/B vssd1 vssd1 vccd1 vccd1 _17899_/A sky130_fd_sc_hd__and2_1
X_19637_ _19638_/CLK _19637_/D vssd1 vssd1 vccd1 vccd1 _19637_/Q sky130_fd_sc_hd__dfxtp_1
X_16849_ _16917_/S vssd1 vssd1 vccd1 vccd1 _16858_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_81_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19568_ _19568_/CLK _19568_/D vssd1 vssd1 vccd1 vccd1 _19568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09321_ _18979_/Q vssd1 vssd1 vccd1 vccd1 _11056_/A sky130_fd_sc_hd__clkbuf_2
X_18519_ _18519_/CLK _18519_/D vssd1 vssd1 vccd1 vccd1 _18519_/Q sky130_fd_sc_hd__dfxtp_2
X_19499_ _19791_/CLK _19499_/D vssd1 vssd1 vccd1 vccd1 _19499_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17725__A2 _13334_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _18573_/Q _18572_/Q _18571_/Q _18570_/Q vssd1 vssd1 vccd1 vccd1 _11519_/A
+ sky130_fd_sc_hd__or4_4
XANTENNA__14539__A2 _12763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09183_ _10379_/A vssd1 vssd1 vccd1 vccd1 _09184_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__18206__A _19856_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14671__A1_N input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12722__A1 _19671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17256__S _17258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_33_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12701__B _18630_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17780__A _17780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09577__S1 _10331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10860_ _18591_/Q _19280_/Q _10860_/S vssd1 vssd1 vccd1 vccd1 _10860_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09519_ _09315_/A _09485_/Y _09503_/X _09506_/Y _09518_/Y vssd1 vssd1 vccd1 vccd1
+ _09519_/X sky130_fd_sc_hd__o32a_1
XFILLER_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13532__B _13536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10648__S _10648_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10791_ _10791_/A vssd1 vssd1 vccd1 vccd1 _10899_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _12530_/A _12686_/A _12791_/A vssd1 vssd1 vccd1 vccd1 _12622_/B sky130_fd_sc_hd__or3_2
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12461_ _12461_/A vssd1 vssd1 vccd1 vccd1 _12461_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14200_ _14297_/A _14203_/A vssd1 vssd1 vccd1 vccd1 _14200_/X sky130_fd_sc_hd__or2_1
X_11412_ _11412_/A vssd1 vssd1 vccd1 vccd1 _12519_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15180_ _15180_/A vssd1 vssd1 vccd1 vccd1 _18663_/D sky130_fd_sc_hd__clkbuf_1
X_12392_ _13388_/A _12393_/C _18378_/Q vssd1 vssd1 vccd1 vccd1 _12392_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_153_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14131_ _13821_/A _14172_/B _14130_/Y _13594_/X vssd1 vssd1 vccd1 vccd1 _14131_/Y
+ sky130_fd_sc_hd__o211ai_1
X_11343_ _11346_/A _11343_/B _11343_/C vssd1 vssd1 vccd1 vccd1 _11343_/X sky130_fd_sc_hd__and3b_2
XFILLER_165_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12164__A _19747_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14062_ _14142_/A _14062_/B vssd1 vssd1 vccd1 vccd1 _14062_/X sky130_fd_sc_hd__or2_1
X_11274_ _11267_/X _11274_/B _11274_/C _11274_/D vssd1 vssd1 vccd1 vccd1 _11274_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_4_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13013_ _13015_/A _13015_/C _13012_/Y vssd1 vssd1 vccd1 vccd1 _18316_/D sky130_fd_sc_hd__o21a_1
XANTENNA__12713__B2 _18630_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10225_ _18834_/Q _19388_/Q _19550_/Q _18802_/Q _10224_/X _09486_/X vssd1 vssd1 vccd1
+ vccd1 _10226_/B sky130_fd_sc_hd__mux4_1
X_18870_ _19003_/CLK _18870_/D vssd1 vssd1 vccd1 vccd1 _18870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17652__A1 _17651_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17821_ _15191_/X _19712_/Q _17827_/S vssd1 vssd1 vccd1 vccd1 _17822_/A sky130_fd_sc_hd__mux2_1
X_10156_ _09984_/X _10153_/X _10155_/X vssd1 vssd1 vccd1 vccd1 _10156_/X sky130_fd_sc_hd__a21o_1
XFILLER_95_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17752_ _17751_/A _17751_/C _15027_/A vssd1 vssd1 vccd1 vccd1 _17752_/Y sky130_fd_sc_hd__o21ai_1
X_14964_ _16813_/A vssd1 vssd1 vccd1 vccd1 _14964_/X sky130_fd_sc_hd__clkbuf_2
X_10087_ _10167_/A vssd1 vssd1 vccd1 vccd1 _10120_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10412__A _10412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16703_ _19294_/Q _16702_/X _16703_/S vssd1 vssd1 vccd1 vccd1 _16704_/A sky130_fd_sc_hd__mux2_1
X_13915_ _13913_/X _13914_/X _14121_/S vssd1 vssd1 vccd1 vccd1 _13915_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17683_ _17683_/A _18473_/Q _17683_/C vssd1 vssd1 vccd1 vccd1 _17691_/B sky130_fd_sc_hd__or3_1
X_14895_ _14883_/A _14894_/C _18474_/Q vssd1 vssd1 vccd1 vccd1 _14896_/C sky130_fd_sc_hd__a21oi_1
XFILLER_75_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19422_ _19616_/CLK _19422_/D vssd1 vssd1 vccd1 vccd1 _19422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16634_ _16634_/A vssd1 vssd1 vccd1 vccd1 _19272_/D sky130_fd_sc_hd__clkbuf_1
X_13846_ _13846_/A vssd1 vssd1 vccd1 vccd1 _13846_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19353_ _19708_/CLK _19353_/D vssd1 vssd1 vccd1 vccd1 _19353_/Q sky130_fd_sc_hd__dfxtp_1
X_13777_ _13773_/X _13776_/X _13968_/S vssd1 vssd1 vccd1 vccd1 _13777_/X sky130_fd_sc_hd__mux2_1
X_16565_ _19238_/Q _15577_/X _16569_/S vssd1 vssd1 vccd1 vccd1 _16566_/A sky130_fd_sc_hd__mux2_1
X_10989_ _10992_/A _10986_/X _10988_/X vssd1 vssd1 vccd1 vccd1 _10989_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18304_ _19790_/CLK _18304_/D vssd1 vssd1 vccd1 vccd1 _18304_/Q sky130_fd_sc_hd__dfxtp_1
X_15516_ _16771_/A vssd1 vssd1 vccd1 vccd1 _15516_/X sky130_fd_sc_hd__clkbuf_2
X_12728_ _13106_/B _12714_/X _12727_/X _13516_/B _12765_/A vssd1 vssd1 vccd1 vccd1
+ _12728_/X sky130_fd_sc_hd__o32a_1
X_19284_ _19726_/CLK _19284_/D vssd1 vssd1 vccd1 vccd1 _19284_/Q sky130_fd_sc_hd__dfxtp_1
X_16496_ _16496_/A vssd1 vssd1 vccd1 vccd1 _19207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18235_ _18250_/A _18239_/C vssd1 vssd1 vccd1 vccd1 _18235_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12659_ _14648_/A vssd1 vssd1 vccd1 vccd1 _12660_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15447_ _15447_/A vssd1 vssd1 vccd1 vccd1 _18766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18166_ _18199_/A vssd1 vssd1 vccd1 vccd1 _18197_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11897__B _13614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15378_ _18737_/Q _15191_/X _15384_/S vssd1 vssd1 vccd1 vccd1 _15379_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17117_ _16819_/X _19458_/Q _17119_/S vssd1 vssd1 vccd1 vccd1 _17118_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17865__A _18225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14329_ _13784_/X _14327_/X _14328_/Y _15123_/A vssd1 vssd1 vccd1 vccd1 _14329_/X
+ sky130_fd_sc_hd__a31o_1
X_18097_ _18097_/A vssd1 vssd1 vccd1 vccd1 _18102_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17048_ _17048_/A vssd1 vssd1 vccd1 vccd1 _19427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09870_ _19268_/Q _19039_/Q _18970_/Q _19364_/Q _09866_/X _09869_/X vssd1 vssd1 vccd1
+ vccd1 _09871_/B sky130_fd_sc_hd__mux4_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11063__S0 _10932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12802__A _18173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10191__A1 _10177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18999_ _19642_/CLK _18999_/D vssd1 vssd1 vccd1 vccd1 _18999_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14457__A1 _11984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11137__B _12486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09884__A1 _09320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11691__A1 _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11118__S1 _10390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16944__A _16990_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11153__A _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09304_ _09624_/A _09624_/B vssd1 vssd1 vccd1 vccd1 _09305_/A sky130_fd_sc_hd__and2_2
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09235_ _09856_/A _09235_/B vssd1 vssd1 vccd1 vccd1 _09235_/X sky130_fd_sc_hd__or2_1
XFILLER_142_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09166_ _19692_/Q vssd1 vssd1 vccd1 vccd1 _10910_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09558__A _10348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09097_ _11320_/A vssd1 vssd1 vccd1 vccd1 _11534_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11054__S0 _10932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12712__A _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10010_ _18607_/Q _19296_/Q _10010_/S vssd1 vssd1 vccd1 vccd1 _10010_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09999_ _19619_/Q _19457_/Q _18903_/Q _18673_/Q _09976_/A _09763_/A vssd1 vssd1 vccd1
+ vccd1 _09999_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14448__A1 _11849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11328__A _11513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11961_ _18360_/Q _13246_/A _11962_/D _18361_/Q vssd1 vssd1 vccd1 vccd1 _11961_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__17398__A0 _16752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14639__A _14673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10912_ _10906_/X _10908_/X _10911_/X _10928_/A _10827_/A vssd1 vssd1 vccd1 vccd1
+ _10917_/B sky130_fd_sc_hd__o221a_1
X_13700_ _13711_/B vssd1 vssd1 vccd1 vccd1 _14150_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14680_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14680_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11892_ _12474_/B _11831_/X _12023_/B _11513_/A vssd1 vssd1 vccd1 vccd1 _14045_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13631_ _13936_/B _12355_/A _13657_/S vssd1 vssd1 vccd1 vccd1 _13631_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10843_ _18758_/Q _18987_/Q _18918_/Q _19216_/Q _11050_/S _10785_/A vssd1 vssd1 vccd1
+ vccd1 _10844_/B sky130_fd_sc_hd__mux4_1
XFILLER_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09627__A1 _09430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16350_ _16350_/A vssd1 vssd1 vccd1 vccd1 _19143_/D sky130_fd_sc_hd__clkbuf_1
X_13562_ _13570_/A _13536_/A _13537_/A _18425_/Q vssd1 vssd1 vccd1 vccd1 _13563_/B
+ sky130_fd_sc_hd__a22o_1
X_10774_ _10774_/A vssd1 vssd1 vccd1 vccd1 _10774_/X sky130_fd_sc_hd__buf_2
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12513_ _12766_/A vssd1 vssd1 vccd1 vccd1 _13171_/A sky130_fd_sc_hd__clkbuf_4
X_15301_ _15301_/A vssd1 vssd1 vccd1 vccd1 _18703_/D sky130_fd_sc_hd__clkbuf_1
X_16281_ _16131_/X _19113_/Q _16283_/S vssd1 vssd1 vccd1 vccd1 _16282_/A sky130_fd_sc_hd__mux2_1
X_13493_ _18405_/Q _13346_/X _13497_/S vssd1 vssd1 vccd1 vccd1 _13494_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16065__S _16065_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18020_ _18207_/A _18023_/A vssd1 vssd1 vccd1 vccd1 _19792_/D sky130_fd_sc_hd__nor2_1
XFILLER_145_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12444_ _11205_/A _18521_/Q _12444_/S vssd1 vssd1 vccd1 vccd1 _12446_/B sky130_fd_sc_hd__mux2_8
X_15232_ _16734_/A vssd1 vssd1 vccd1 vccd1 _15232_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15163_ _18658_/Q _15162_/X _15169_/S vssd1 vssd1 vccd1 vccd1 _15164_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11510__B _14568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17322__A0 _16743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12375_ _12290_/B _12313_/A _12371_/X _12374_/X vssd1 vssd1 vccd1 vccd1 _12385_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_154_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14114_ _14037_/X _14106_/X _14113_/Y _13594_/A vssd1 vssd1 vccd1 vccd1 _14114_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11326_ _18583_/Q vssd1 vssd1 vccd1 vccd1 _11513_/A sky130_fd_sc_hd__buf_2
X_15094_ _15094_/A vssd1 vssd1 vccd1 vccd1 _18623_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14687__A1 _11517_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14687__B2 input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18922_ _19444_/CLK _18922_/D vssd1 vssd1 vccd1 vccd1 _18922_/Q sky130_fd_sc_hd__dfxtp_1
X_14045_ _14045_/A _14045_/B vssd1 vssd1 vccd1 vccd1 _14045_/Y sky130_fd_sc_hd__nor2_1
X_11257_ _11257_/A _11257_/B vssd1 vssd1 vccd1 vccd1 _11258_/C sky130_fd_sc_hd__or2_1
XANTENNA__09789__S1 _09841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12622__A _14562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12698__B1 _18205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10208_ _09215_/A _10199_/X _10203_/X _10207_/X _09134_/A vssd1 vssd1 vccd1 vccd1
+ _10208_/X sky130_fd_sc_hd__a311o_1
XFILLER_95_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18853_ _18853_/CLK _18853_/D vssd1 vssd1 vccd1 vccd1 _18853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11188_ _18614_/Q _19303_/Q _11188_/S vssd1 vssd1 vccd1 vccd1 _11189_/B sky130_fd_sc_hd__mux2_1
XFILLER_68_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14439__A1 _19730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17624__S _17628_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17804_ _17804_/A vssd1 vssd1 vccd1 vccd1 _19704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10139_ _19520_/Q _19134_/Q _19584_/Q _18740_/Q _10125_/X _09867_/A vssd1 vssd1 vccd1
+ vccd1 _10140_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15100__A2 _13566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18784_ _19727_/CLK _18784_/D vssd1 vssd1 vccd1 vccd1 _18784_/Q sky130_fd_sc_hd__dfxtp_1
X_15996_ _16018_/A vssd1 vssd1 vccd1 vccd1 _16005_/S sky130_fd_sc_hd__buf_4
X_17735_ _19682_/Q _17734_/X _17772_/S vssd1 vssd1 vccd1 vccd1 _17736_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11122__A0 _18830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14947_ _18446_/Q _15018_/A _14946_/X _14980_/A vssd1 vssd1 vccd1 vccd1 _14947_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15144__S _15153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17666_ _17666_/A vssd1 vssd1 vccd1 vccd1 _19670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12870__B1 _12869_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09961__S1 _09936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14878_ _16686_/A vssd1 vssd1 vccd1 vccd1 _16790_/A sky130_fd_sc_hd__buf_2
XFILLER_36_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19405_ _19631_/CLK _19405_/D vssd1 vssd1 vccd1 vccd1 _19405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16617_ _19264_/Q vssd1 vssd1 vccd1 vccd1 _16618_/A sky130_fd_sc_hd__clkbuf_1
X_13829_ _11624_/Y _13827_/X _13828_/X vssd1 vssd1 vccd1 vccd1 _13829_/X sky130_fd_sc_hd__a21o_1
XFILLER_63_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13414__A2 _13412_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17597_ _19656_/Q _16832_/A _17601_/S vssd1 vssd1 vccd1 vccd1 _17598_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19336_ _19626_/CLK _19336_/D vssd1 vssd1 vccd1 vccd1 _19336_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09713__S1 _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16548_ _16548_/A vssd1 vssd1 vccd1 vccd1 _19230_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19267_ _19589_/CLK _19267_/D vssd1 vssd1 vccd1 vccd1 _19267_/Q sky130_fd_sc_hd__dfxtp_1
X_16479_ _16479_/A vssd1 vssd1 vccd1 vccd1 _19199_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14284__A _14284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18218_ _19860_/Q _18215_/B _18217_/Y vssd1 vssd1 vccd1 vccd1 _19860_/D sky130_fd_sc_hd__o21a_1
XANTENNA__09378__A _10593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19198_ _19660_/CLK _19198_/D vssd1 vssd1 vccd1 vccd1 _19198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18149_ _18165_/A _18149_/B _18150_/B vssd1 vssd1 vccd1 vccd1 _19836_/D sky130_fd_sc_hd__nor3_1
XANTENNA__16703__S _16703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09922_ _09217_/X _09917_/X _09919_/X _09921_/X _09854_/A vssd1 vssd1 vccd1 vccd1
+ _09922_/X sky130_fd_sc_hd__a221o_2
XFILLER_116_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11036__S0 _10959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13628__A _13650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09853_ _09905_/A _09850_/X _09852_/X _09231_/X vssd1 vssd1 vccd1 vccd1 _09854_/C
+ sky130_fd_sc_hd__o211a_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11148__A _11148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09784_ _19427_/Q _19203_/Q _19720_/Q _19171_/Q _09782_/X _09783_/X vssd1 vssd1 vccd1
+ vccd1 _09784_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09841__A _09841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12684__B1_N _12600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14850__A1 _12726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14178__B _14178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16674__A _16741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13169__A1 _13112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09218_ _09165_/X _09189_/X _09191_/X _09856_/A _09217_/X vssd1 vssd1 vccd1 vccd1
+ _09233_/B sky130_fd_sc_hd__o221a_1
XFILLER_167_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09288__A _18533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10490_ _19414_/Q _19190_/Q _19707_/Q _19158_/Q _10450_/S _09587_/A vssd1 vssd1 vccd1
+ vccd1 _10490_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12426__B _14324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09149_ _09149_/A vssd1 vssd1 vccd1 vccd1 _09165_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14118__A0 _18439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12160_ _12160_/A _13598_/A vssd1 vssd1 vccd1 vccd1 _12161_/B sky130_fd_sc_hd__nor2_1
XFILLER_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11111_ _11111_/A _11110_/X vssd1 vssd1 vccd1 vccd1 _11111_/X sky130_fd_sc_hd__or2b_1
XANTENNA_clkbuf_2_2_0_clock_A clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12091_ _12091_/A vssd1 vssd1 vccd1 vccd1 _17711_/A sky130_fd_sc_hd__buf_4
XFILLER_123_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11984__C _17878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11042_ _18817_/Q _19371_/Q _19533_/Q _18785_/Q _10919_/X _10920_/X vssd1 vssd1 vccd1
+ vccd1 _11042_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10155__A1 _09173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16849__A _16917_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17444__S _17446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15850_ _14929_/X _18931_/Q _15852_/S vssd1 vssd1 vccd1 vccd1 _15851_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09751__A _18452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14801_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14801_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_input20_A io_dbus_rdata[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _15781_/A vssd1 vssd1 vccd1 vccd1 _18900_/D sky130_fd_sc_hd__clkbuf_1
X_12993_ _12993_/A _18311_/Q _12993_/C vssd1 vssd1 vccd1 vccd1 _12994_/C sky130_fd_sc_hd__and3_1
X_17520_ _17520_/A vssd1 vssd1 vccd1 vccd1 _17529_/S sky130_fd_sc_hd__buf_4
XFILLER_18_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14732_ _14842_/A vssd1 vssd1 vccd1 vccd1 _14732_/X sky130_fd_sc_hd__buf_2
XANTENNA__09943__S1 _09869_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11944_ _13524_/B _12024_/A _11943_/X vssd1 vssd1 vccd1 vccd1 _11944_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_91_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _16829_/X _19591_/Q _17457_/S vssd1 vssd1 vccd1 vccd1 _17452_/A sky130_fd_sc_hd__mux2_1
X_11875_ _11810_/A _11843_/A _11842_/A _13658_/A vssd1 vssd1 vccd1 vccd1 _11875_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14663_ input46/X _14640_/X _14643_/X _13524_/B vssd1 vssd1 vccd1 vccd1 _15952_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output107_A _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _19166_/Q _15551_/X _16402_/S vssd1 vssd1 vccd1 vccd1 _16403_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10826_ _19633_/Q _19050_/Q _19087_/Q _18693_/Q _09152_/A _10740_/A vssd1 vssd1 vccd1
+ vccd1 _10826_/X sky130_fd_sc_hd__mux4_2
X_13614_ _13614_/A vssd1 vssd1 vccd1 vccd1 _14045_/B sky130_fd_sc_hd__buf_2
XFILLER_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17382_ _17382_/A vssd1 vssd1 vccd1 vccd1 _19560_/D sky130_fd_sc_hd__clkbuf_1
X_14594_ input34/X vssd1 vssd1 vccd1 vccd1 _14594_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_2_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19121_ _19635_/CLK _19121_/D vssd1 vssd1 vccd1 vccd1 _19121_/Q sky130_fd_sc_hd__dfxtp_1
X_16333_ _16333_/A vssd1 vssd1 vccd1 vccd1 _19135_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13720__B _13720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10757_ _09210_/A _10750_/X _10752_/X _10756_/X _09245_/A vssd1 vssd1 vccd1 vccd1
+ _10757_/X sky130_fd_sc_hd__a311o_2
X_13545_ _13578_/A _13545_/B _13545_/C vssd1 vssd1 vccd1 vccd1 _13545_/X sky130_fd_sc_hd__and3b_1
XANTENNA_clkbuf_leaf_155_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10091__B1 _10007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11521__A _11561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09198__A _11097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19052_ _19635_/CLK _19052_/D vssd1 vssd1 vccd1 vccd1 _19052_/Q sky130_fd_sc_hd__dfxtp_1
X_16264_ _16106_/X _19105_/Q _16268_/S vssd1 vssd1 vccd1 vccd1 _16265_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13476_ _13476_/A vssd1 vssd1 vccd1 vccd1 _18397_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10630__A2 _10620_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10688_ _18824_/Q _19378_/Q _19540_/Q _18792_/Q _10669_/A _10670_/X vssd1 vssd1 vccd1
+ vccd1 _10688_/X sky130_fd_sc_hd__mux4_2
XFILLER_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18003_ _19786_/Q _18006_/C _17993_/X vssd1 vssd1 vccd1 vccd1 _18003_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_173_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15215_ _15215_/A vssd1 vssd1 vccd1 vccd1 _18674_/D sky130_fd_sc_hd__clkbuf_1
X_12427_ _12427_/A _12426_/X vssd1 vssd1 vccd1 vccd1 _12431_/A sky130_fd_sc_hd__or2b_2
X_16195_ _16195_/A vssd1 vssd1 vccd1 vccd1 _19070_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14832__A _16673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15146_ _16648_/A vssd1 vssd1 vccd1 vccd1 _15146_/X sky130_fd_sc_hd__clkbuf_2
X_12358_ _14284_/A vssd1 vssd1 vccd1 vccd1 _12358_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11309_ _11736_/A vssd1 vssd1 vccd1 vccd1 _11692_/A sky130_fd_sc_hd__clkbuf_2
X_15077_ _15076_/X _18617_/Q _15077_/S vssd1 vssd1 vccd1 vccd1 _15078_/A sky130_fd_sc_hd__mux2_1
X_12289_ _12240_/A _12240_/B _12265_/A _12288_/Y vssd1 vssd1 vccd1 vccd1 _12290_/B
+ sky130_fd_sc_hd__a31o_2
XANTENNA__13332__A1 _19845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18905_ _19720_/CLK _18905_/D vssd1 vssd1 vccd1 vccd1 _18905_/Q sky130_fd_sc_hd__dfxtp_1
X_14028_ _14023_/Y _14025_/Y _14027_/X vssd1 vssd1 vccd1 vccd1 _14028_/X sky130_fd_sc_hd__a21o_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18836_ _19584_/CLK _18836_/D vssd1 vssd1 vccd1 vccd1 _18836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11894__A1 _12057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18767_ _19223_/CLK _18767_/D vssd1 vssd1 vccd1 vccd1 _18767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15979_ _14792_/X _18989_/Q _15983_/S vssd1 vssd1 vccd1 vccd1 _15980_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17718_ _19679_/Q _17717_/X _17718_/S vssd1 vssd1 vccd1 vccd1 _17719_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09934__S1 _09869_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18698_ _19638_/CLK _18698_/D vssd1 vssd1 vccd1 vccd1 _18698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17649_ _18466_/Q _18467_/Q _17649_/C vssd1 vssd1 vccd1 vccd1 _17656_/B sky130_fd_sc_hd__or3_1
XFILLER_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13333__D _14958_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19319_ _19513_/CLK _19319_/D vssd1 vssd1 vccd1 vccd1 _19319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17529__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15848__A0 _14918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09870__S0 _09866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11009__S0 _18977_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13323__A1 _12656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09905_ _09905_/A _09905_/B vssd1 vssd1 vccd1 vccd1 _09905_/X sky130_fd_sc_hd__or2_1
XFILLER_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09836_ _09819_/A _09831_/X _09835_/X vssd1 vssd1 vccd1 vccd1 _09836_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_101_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10232__S1 _11111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ _10115_/A _09767_/B vssd1 vssd1 vccd1 vccd1 _09767_/X sky130_fd_sc_hd__and2_1
XFILLER_58_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _11157_/S vssd1 vssd1 vccd1 vccd1 _10256_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_55_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11325__B _14575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14917__A _16696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ _12072_/A vssd1 vssd1 vccd1 vccd1 _17221_/A sky130_fd_sc_hd__buf_2
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _19411_/Q _19187_/Q _19704_/Q _19155_/Q _10353_/A _10548_/X vssd1 vssd1 vccd1
+ vccd1 _10611_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11591_ _10857_/X _11035_/X _11044_/X _11046_/Y vssd1 vssd1 vccd1 vccd1 _11591_/Y
+ sky130_fd_sc_hd__o31ai_4
XFILLER_22_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13330_ _18256_/Q _12651_/X _12753_/X _19781_/Q vssd1 vssd1 vccd1 vccd1 _14958_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10542_ _09170_/A _10541_/X _09451_/A vssd1 vssd1 vccd1 vccd1 _10542_/X sky130_fd_sc_hd__a21o_1
XFILLER_167_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13261_ _18360_/Q _13295_/B vssd1 vssd1 vccd1 vccd1 _13261_/X sky130_fd_sc_hd__or2_1
X_10473_ _09212_/A _10464_/X _10468_/X _10472_/X _10373_/A vssd1 vssd1 vccd1 vccd1
+ _10473_/X sky130_fd_sc_hd__a311o_4
XANTENNA__16343__S _16351_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12212_ _12235_/A _12212_/B vssd1 vssd1 vccd1 vccd1 _14211_/A sky130_fd_sc_hd__xnor2_4
X_15000_ _15000_/A vssd1 vssd1 vccd1 vccd1 _15000_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13562__A1 _13570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13192_ _19829_/Q vssd1 vssd1 vccd1 vccd1 _18131_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_163_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input68_A io_irq_m2_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12143_ _19745_/Q _12144_/C _19746_/Q vssd1 vssd1 vccd1 vccd1 _12145_/A sky130_fd_sc_hd__a21oi_1
XFILLER_135_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14802__D input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09518__B1 _09681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12074_ _13295_/A _12075_/C _18365_/Q vssd1 vssd1 vccd1 vccd1 _12074_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16951_ _16787_/X _19384_/Q _16953_/S vssd1 vssd1 vccd1 vccd1 _16952_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11025_ _19243_/Q _19014_/Q _18945_/Q _19339_/Q _10919_/X _10920_/X vssd1 vssd1 vccd1
+ vccd1 _11026_/B sky130_fd_sc_hd__mux4_2
X_15902_ _14821_/X _18954_/Q _15902_/S vssd1 vssd1 vccd1 vccd1 _15903_/A sky130_fd_sc_hd__mux2_1
X_19670_ _19687_/CLK _19670_/D vssd1 vssd1 vccd1 vccd1 _19670_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_49_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16882_ _16904_/A vssd1 vssd1 vccd1 vccd1 _16891_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_38_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_6_0_clock_A clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_81_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09481__A _09481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18621_ _18623_/CLK _18621_/D vssd1 vssd1 vccd1 vccd1 _18621_/Q sky130_fd_sc_hd__dfxtp_2
X_15833_ _14833_/X _18923_/Q _15841_/S vssd1 vssd1 vccd1 vccd1 _15834_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14814__A1 _18435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18552_ _19481_/CLK _18552_/D vssd1 vssd1 vccd1 vccd1 _18552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09916__S1 _09783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15764_ _15764_/A vssd1 vssd1 vccd1 vccd1 _18892_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _12997_/A _12982_/C vssd1 vssd1 vccd1 vccd1 _12976_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09297__A2 _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17503_ _19614_/Q _16696_/X _17507_/S vssd1 vssd1 vccd1 vccd1 _17504_/A sky130_fd_sc_hd__mux2_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _18533_/Q vssd1 vssd1 vccd1 vccd1 _16919_/A sky130_fd_sc_hd__clkbuf_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _19738_/Q vssd1 vssd1 vccd1 vccd1 _11984_/A sky130_fd_sc_hd__buf_4
X_18483_ _18519_/CLK _18483_/D vssd1 vssd1 vccd1 vccd1 _18483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15695_ _18862_/Q _15532_/X _15697_/S vssd1 vssd1 vccd1 vccd1 _15696_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14027__C1 _13711_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15422__S _15426_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17434_ _17434_/A vssd1 vssd1 vccd1 vccd1 _19583_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14646_ input40/X _14640_/X _14643_/X _14551_/A vssd1 vssd1 vccd1 vccd1 _17774_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_11858_ _13215_/A _11758_/X _11888_/D _11994_/A vssd1 vssd1 vccd1 vccd1 _11858_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__14042__A2 _14045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12053__A1 _12067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17365_ _17376_/A vssd1 vssd1 vccd1 vccd1 _17374_/S sky130_fd_sc_hd__buf_4
X_10809_ _09408_/A _10801_/X _10803_/X _10808_/X _09391_/A vssd1 vssd1 vccd1 vccd1
+ _10809_/X sky130_fd_sc_hd__a311o_2
X_11789_ _11994_/A vssd1 vssd1 vccd1 vccd1 _11790_/A sky130_fd_sc_hd__clkbuf_2
X_14577_ _14577_/A vssd1 vssd1 vccd1 vccd1 _14577_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19104_ _19812_/CLK _19104_/D vssd1 vssd1 vccd1 vccd1 _19104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16316_ _16077_/X _19128_/Q _16318_/S vssd1 vssd1 vccd1 vccd1 _16317_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13528_ _11628_/C _13524_/X _13545_/C _13545_/B _13527_/X vssd1 vssd1 vccd1 vccd1
+ _13529_/D sky130_fd_sc_hd__o2111a_1
X_17296_ _19522_/Q _16709_/X _17302_/S vssd1 vssd1 vccd1 vccd1 _17297_/A sky130_fd_sc_hd__mux2_1
X_19035_ _19818_/CLK _19035_/D vssd1 vssd1 vccd1 vccd1 _19035_/Q sky130_fd_sc_hd__dfxtp_1
X_16247_ _16247_/A vssd1 vssd1 vccd1 vccd1 _19097_/D sky130_fd_sc_hd__clkbuf_1
X_13459_ _13459_/A vssd1 vssd1 vccd1 vccd1 _18389_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14562__A _14562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16253__S _16257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13553__A1 _09109_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput104 _11899_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[9] sky130_fd_sc_hd__buf_2
XANTENNA__14750__B1 _14749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput115 _12481_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[13] sky130_fd_sc_hd__buf_2
X_16178_ _16178_/A vssd1 vssd1 vccd1 vccd1 _19062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput126 _12496_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[23] sky130_fd_sc_hd__buf_2
Xoutput137 _12465_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[4] sky130_fd_sc_hd__buf_2
Xoutput148 _17880_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[13] sky130_fd_sc_hd__buf_2
XFILLER_126_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15129_ _18647_/Q _15123_/X _15125_/X _11199_/A vssd1 vssd1 vccd1 vccd1 _18647_/D
+ sky130_fd_sc_hd__a22o_1
Xoutput159 _17900_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[23] sky130_fd_sc_hd__buf_2
XFILLER_142_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19868_ _19871_/CLK _19868_/D vssd1 vssd1 vccd1 vccd1 _19868_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10214__S1 _09697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12810__A _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09391__A _09391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09621_ _09621_/A vssd1 vssd1 vccd1 vccd1 _09621_/X sky130_fd_sc_hd__buf_2
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18819_ _19537_/CLK _18819_/D vssd1 vssd1 vccd1 vccd1 _18819_/Q sky130_fd_sc_hd__dfxtp_1
X_19799_ _19804_/CLK _19799_/D vssd1 vssd1 vccd1 vccd1 _19799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14805__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15488__C_N _16919_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17812__S _17816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ _10309_/A vssd1 vssd1 vccd1 vccd1 _09772_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09907__S1 _09783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09483_ _09662_/A vssd1 vssd1 vccd1 vccd1 _09483_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__16428__S _16428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14737__A _14737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09566__A _10313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13088__A _13088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17783__A _17783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10453__S1 _11111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_103_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10205__S1 _10080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09819_ _09819_/A _09819_/B vssd1 vssd1 vccd1 vccd1 _09819_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11981__D _19739_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12830_ _18259_/Q _12830_/B _12830_/C vssd1 vssd1 vccd1 vccd1 _12831_/C sky130_fd_sc_hd__and3_1
XFILLER_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _14516_/S vssd1 vssd1 vccd1 vccd1 _14565_/A sky130_fd_sc_hd__buf_2
XANTENNA__16338__S _16340_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09684__C1 _09394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10294__B1 _09681_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14500_ _18520_/Q _19758_/Q _14502_/S vssd1 vssd1 vccd1 vccd1 _14501_/A sky130_fd_sc_hd__mux2_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _12072_/A vssd1 vssd1 vccd1 vccd1 _12696_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _15480_/A vssd1 vssd1 vccd1 vccd1 _18781_/D sky130_fd_sc_hd__clkbuf_1
X_12692_ _14577_/A vssd1 vssd1 vccd1 vccd1 _12692_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_15_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _13584_/B _13570_/D _11643_/C _13571_/B vssd1 vssd1 vccd1 vccd1 _11645_/B
+ sky130_fd_sc_hd__or4b_1
X_14431_ _14431_/A _14431_/B _14431_/C _13529_/A vssd1 vssd1 vccd1 vccd1 _14432_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_30_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17150_ _18429_/Q _17628_/S _17149_/Y vssd1 vssd1 vccd1 vccd1 _17150_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_opt_1_0_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
X_14362_ _14362_/A vssd1 vssd1 vccd1 vccd1 _18465_/D sky130_fd_sc_hd__clkbuf_1
X_11574_ _11735_/S vssd1 vssd1 vccd1 vccd1 _15095_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_28_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10141__S0 _09734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput17 io_dbus_rdata[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_2
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16101_ _16099_/X _19034_/Q _16113_/S vssd1 vssd1 vccd1 vccd1 _16102_/A sky130_fd_sc_hd__mux2_1
Xinput28 io_dbus_rdata[5] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13313_ _12559_/X _13311_/X _13312_/X _13282_/X vssd1 vssd1 vccd1 vccd1 _18366_/D
+ sky130_fd_sc_hd__o211a_1
Xinput39 io_ibus_inst[14] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10525_ _18827_/Q _19381_/Q _19543_/Q _18795_/Q _10387_/S _10501_/X vssd1 vssd1 vccd1
+ vccd1 _10525_/X sky130_fd_sc_hd__mux4_2
XFILLER_128_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14293_ _14328_/A _14293_/B vssd1 vssd1 vccd1 vccd1 _14293_/Y sky130_fd_sc_hd__nand2_1
X_17081_ _17081_/A vssd1 vssd1 vccd1 vccd1 _19441_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14813__C _14813_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13244_ _18628_/Q _14813_/B _14813_/C _14813_/D vssd1 vssd1 vccd1 vccd1 _13244_/X
+ sky130_fd_sc_hd__or4_1
X_16032_ _16032_/A vssd1 vssd1 vccd1 vccd1 _19013_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09739__B1 _09317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10456_ _10442_/A _10453_/X _10455_/X vssd1 vssd1 vccd1 vccd1 _10456_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09834__S0 _09874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17693__A _17693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13175_ _19473_/Q _12741_/X _13173_/X _13174_/X vssd1 vssd1 vccd1 vccd1 _13175_/X
+ sky130_fd_sc_hd__a211o_1
X_10387_ _18863_/Q _19321_/Q _10387_/S vssd1 vssd1 vccd1 vccd1 _10388_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16801__S _16807_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12126_ _12126_/A vssd1 vssd1 vccd1 vccd1 _12226_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17983_ _19779_/Q _17981_/B _17982_/Y vssd1 vssd1 vccd1 vccd1 _19779_/D sky130_fd_sc_hd__o21a_1
XFILLER_97_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19722_ _19722_/CLK _19722_/D vssd1 vssd1 vccd1 vccd1 _19722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16934_ _16761_/X _19376_/Q _16942_/S vssd1 vssd1 vccd1 vccd1 _16935_/A sky130_fd_sc_hd__mux2_1
X_12057_ _12057_/A vssd1 vssd1 vccd1 vccd1 _12348_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11008_ _19404_/Q _19180_/Q _19697_/Q _19148_/Q _09336_/A _10940_/X vssd1 vssd1 vccd1
+ vccd1 _11008_/X sky130_fd_sc_hd__mux4_2
XFILLER_78_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19653_ _19718_/CLK _19653_/D vssd1 vssd1 vccd1 vccd1 _19653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16865_ _19346_/Q _16664_/X _16869_/S vssd1 vssd1 vccd1 vccd1 _16866_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18604_ _19584_/CLK _18604_/D vssd1 vssd1 vccd1 vccd1 _18604_/Q sky130_fd_sc_hd__dfxtp_1
X_15816_ _15816_/A vssd1 vssd1 vccd1 vccd1 _18915_/D sky130_fd_sc_hd__clkbuf_1
X_19584_ _19584_/CLK _19584_/D vssd1 vssd1 vccd1 vccd1 _19584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10150__A _11139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16796_ _16796_/A vssd1 vssd1 vccd1 vccd1 _19322_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14263__A2 _14265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18535_ _18567_/CLK _18535_/D vssd1 vssd1 vccd1 vccd1 _18535_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10809__C1 _09391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ _14761_/X _18885_/Q _15747_/S vssd1 vssd1 vccd1 vccd1 _15748_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12959_ _18297_/Q _12959_/B vssd1 vssd1 vccd1 vccd1 _12961_/A sky130_fd_sc_hd__and2_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14557__A _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18466_ _18632_/CLK _18466_/D vssd1 vssd1 vccd1 vccd1 _18466_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15678_ _18854_/Q _15506_/X _15686_/S vssd1 vssd1 vccd1 vccd1 _15679_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10380__S0 _10417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17417_ _17417_/A vssd1 vssd1 vccd1 vccd1 _19575_/D sky130_fd_sc_hd__clkbuf_1
X_14629_ _14629_/A vssd1 vssd1 vccd1 vccd1 _18563_/D sky130_fd_sc_hd__clkbuf_1
X_18397_ _19496_/CLK _18397_/D vssd1 vssd1 vccd1 vccd1 _18397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17348_ _16784_/X _19545_/Q _17352_/S vssd1 vssd1 vccd1 vccd1 _17349_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10588__A1 _10593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17279_ _17279_/A vssd1 vssd1 vccd1 vccd1 _19514_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12805__A _13042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19018_ _19633_/CLK _19018_/D vssd1 vssd1 vccd1 vccd1 _19018_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14723__A0 _14714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15327__S _15333_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10512__A1 _10245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17542__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09604_ _19272_/Q _19043_/Q _18974_/Q _19368_/Q _09734_/A _09610_/A vssd1 vssd1 vccd1
+ vccd1 _09604_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15451__A1 _15187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09535_ _09640_/A vssd1 vssd1 vccd1 vccd1 _10262_/A sky130_fd_sc_hd__buf_2
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14467__A _14591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09466_ _18847_/Q _19401_/Q _19563_/Q _18815_/Q _10465_/S _09142_/A vssd1 vssd1 vccd1
+ vccd1 _09466_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15997__S _16005_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17778__A _17778_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09397_ _18981_/Q vssd1 vssd1 vccd1 vccd1 _10944_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_174_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19726_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10934__S _10934_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10674__S1 _10548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10310_ _10313_/A _10307_/X _10309_/X _09562_/X vssd1 vssd1 vccd1 vccd1 _10310_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09296__A _18574_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11290_ _11565_/A _11565_/B vssd1 vssd1 vccd1 vccd1 _19468_/D sky130_fd_sc_hd__nand2_2
XFILLER_152_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12725__C1 _12724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_189_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19543_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_3_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10241_ _10241_/A vssd1 vssd1 vccd1 vccd1 _10241_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10172_ _19615_/Q _19453_/Q _18899_/Q _18669_/Q _09344_/A _11189_/A vssd1 vssd1 vccd1
+ vccd1 _10173_/B sky130_fd_sc_hd__mux4_1
XFILLER_105_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_112_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19732_/CLK sky130_fd_sc_hd__clkbuf_16
X_14980_ _14980_/A _14980_/B _15002_/C vssd1 vssd1 vccd1 vccd1 _14980_/X sky130_fd_sc_hd__or3_1
XFILLER_94_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13931_ _13931_/A _13931_/B _13931_/C vssd1 vssd1 vccd1 vccd1 _13931_/X sky130_fd_sc_hd__or3_1
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16650_ _16650_/A vssd1 vssd1 vccd1 vccd1 _19277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13862_ _13862_/A _13862_/B _13862_/C vssd1 vssd1 vccd1 vccd1 _13868_/A sky130_fd_sc_hd__or3_1
XFILLER_75_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15601_ _18820_/Q _15500_/X _15603_/S vssd1 vssd1 vccd1 vccd1 _15602_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_127_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _18510_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_170_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12813_ _18254_/Q _18253_/Q _18252_/Q _12813_/D vssd1 vssd1 vccd1 vccd1 _12823_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_16_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16581_ _19246_/Q vssd1 vssd1 vccd1 vccd1 _16582_/A sky130_fd_sc_hd__clkbuf_1
X_13793_ _14003_/A vssd1 vssd1 vccd1 vccd1 _13856_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18320_ _19810_/CLK _18320_/D vssd1 vssd1 vccd1 vccd1 _18320_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13281__A _17892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15532_ _16787_/A vssd1 vssd1 vccd1 vccd1 _15532_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _19492_/Q _12741_/X _12743_/X _18406_/Q vssd1 vssd1 vccd1 vccd1 _12744_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17195__A1 _12559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _19872_/Q _18249_/B _18250_/Y vssd1 vssd1 vccd1 vccd1 _19872_/D sky130_fd_sc_hd__o21a_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _15463_/A vssd1 vssd1 vccd1 vccd1 _18773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _18270_/Q vssd1 vssd1 vccd1 vccd1 _12873_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_31_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17202_ _19487_/Q _17201_/X _17206_/S vssd1 vssd1 vccd1 vccd1 _17203_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15700__S _15708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14414_ _14414_/A vssd1 vssd1 vccd1 vccd1 _18483_/D sky130_fd_sc_hd__clkbuf_1
X_18182_ _19847_/Q _18183_/C _19848_/Q vssd1 vssd1 vccd1 vccd1 _18184_/B sky130_fd_sc_hd__a21oi_1
X_11626_ _15241_/B vssd1 vssd1 vccd1 vccd1 _17611_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15394_ _15394_/A vssd1 vssd1 vccd1 vccd1 _18744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17133_ _17133_/A vssd1 vssd1 vccd1 vccd1 _19465_/D sky130_fd_sc_hd__clkbuf_1
X_14345_ _18460_/Q vssd1 vssd1 vccd1 vccd1 _14743_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11557_ _12469_/B _13532_/A vssd1 vssd1 vccd1 vccd1 _11557_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__13508__A1 _13412_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14705__A0 _11046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17064_ _17463_/A _17064_/B vssd1 vssd1 vccd1 vccd1 _17121_/A sky130_fd_sc_hd__or2_2
X_10508_ _19253_/Q _19024_/Q _18955_/Q _19349_/Q _10387_/S _10501_/X vssd1 vssd1 vccd1
+ vccd1 _10508_/X sky130_fd_sc_hd__mux4_1
X_11488_ _14250_/A vssd1 vssd1 vccd1 vccd1 _14089_/A sky130_fd_sc_hd__clkbuf_4
X_14276_ _14276_/A _14276_/B vssd1 vssd1 vccd1 vccd1 _14276_/X sky130_fd_sc_hd__or2_1
XFILLER_109_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10990__A1 _10821_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16015_ _16015_/A vssd1 vssd1 vccd1 vccd1 _19005_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14181__A1 _14178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13227_ _19800_/Q _12665_/X _12602_/X _18311_/Q _13226_/X vssd1 vssd1 vccd1 vccd1
+ _13228_/B sky130_fd_sc_hd__a221o_2
X_10439_ _19609_/Q _19447_/Q _18893_/Q _18663_/Q _11112_/S _09602_/A vssd1 vssd1 vccd1
+ vccd1 _10440_/B sky130_fd_sc_hd__mux4_1
XFILLER_98_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _18269_/Q _13326_/B _13251_/A _19661_/Q _13157_/X vssd1 vssd1 vccd1 vccd1
+ _13158_/X sky130_fd_sc_hd__a221o_1
XFILLER_69_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15147__S _15153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _11137_/A _18507_/Q _12177_/A vssd1 vssd1 vccd1 vccd1 _13608_/A sky130_fd_sc_hd__mux2_4
X_17966_ _17991_/A _17971_/C vssd1 vssd1 vccd1 vccd1 _17966_/Y sky130_fd_sc_hd__nor2_1
X_13089_ _18335_/Q _11790_/X _12714_/B _13110_/A vssd1 vssd1 vccd1 vccd1 _13089_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12360__A _12361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16917_ _19370_/Q _16740_/X _16917_/S vssd1 vssd1 vccd1 vccd1 _16918_/A sky130_fd_sc_hd__mux2_1
X_19705_ _19726_/CLK _19705_/D vssd1 vssd1 vccd1 vccd1 _19705_/Q sky130_fd_sc_hd__dfxtp_1
X_17897_ _19749_/Q _17886_/X _12224_/Y _14585_/X vssd1 vssd1 vccd1 vccd1 _19749_/D
+ sky130_fd_sc_hd__o211a_1
X_16848_ _16904_/A vssd1 vssd1 vccd1 vccd1 _16917_/S sky130_fd_sc_hd__buf_8
X_19636_ _19636_/CLK _19636_/D vssd1 vssd1 vccd1 vccd1 _19636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15433__A1 _15162_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19567_ _19631_/CLK _19567_/D vssd1 vssd1 vccd1 vccd1 _19567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16779_ _16777_/X _19317_/Q _16791_/S vssd1 vssd1 vccd1 vccd1 _16780_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14287__A _14289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09320_ _09320_/A vssd1 vssd1 vccd1 vccd1 _09320_/X sky130_fd_sc_hd__buf_4
X_18518_ _18519_/CLK _18518_/D vssd1 vssd1 vccd1 vccd1 _18518_/Q sky130_fd_sc_hd__dfxtp_2
X_19498_ _19788_/CLK _19498_/D vssd1 vssd1 vccd1 vccd1 _19498_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_91_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19872_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09251_ _18569_/Q vssd1 vssd1 vccd1 vccd1 _11497_/A sky130_fd_sc_hd__buf_2
XFILLER_167_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18449_ _19634_/CLK _18449_/D vssd1 vssd1 vccd1 vccd1 _18449_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09182_ _11099_/A vssd1 vssd1 vccd1 vccd1 _10379_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10430__B1 _09212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13366__A _18375_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12270__A _19682_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_44_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19722_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_112_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16677__A _16677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17272__S _17280_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15424__A1 _15149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10592__S0 _10511_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09518_ _10498_/A _09516_/X _09681_/A vssd1 vssd1 vccd1 vccd1 _09518_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_59_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19555_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10790_ _10887_/A _10790_/B vssd1 vssd1 vccd1 vccd1 _10790_/X sky130_fd_sc_hd__and2b_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09449_/A vssd1 vssd1 vccd1 vccd1 _10348_/S sky130_fd_sc_hd__clkbuf_4
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14935__A0 _18445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12460_ _12460_/A _12466_/B vssd1 vssd1 vccd1 vccd1 _12461_/A sky130_fd_sc_hd__and2_1
XFILLER_71_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ _12533_/A _12533_/B vssd1 vssd1 vccd1 vccd1 _12540_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12391_ _11706_/X _12389_/X _12390_/X _12072_/X vssd1 vssd1 vccd1 vccd1 _12391_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10664__S _10664_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12445__A _14332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14130_ _14130_/A _14130_/B vssd1 vssd1 vccd1 vccd1 _14130_/Y sky130_fd_sc_hd__nand2_1
X_11342_ _18585_/Q _18560_/Q _11321_/B _18558_/Q vssd1 vssd1 vccd1 vccd1 _11346_/A
+ sky130_fd_sc_hd__or4bb_1
XFILLER_165_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14061_ _14276_/A vssd1 vssd1 vccd1 vccd1 _14142_/A sky130_fd_sc_hd__clkbuf_2
X_11273_ _11225_/B _11145_/A _11272_/Y _11271_/A vssd1 vssd1 vccd1 vccd1 _11274_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16351__S _16351_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input50_A io_ibus_inst[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13012_ _13015_/A _13015_/C _13011_/X vssd1 vssd1 vccd1 vccd1 _13012_/Y sky130_fd_sc_hd__a21oi_1
X_10224_ _10486_/S vssd1 vssd1 vccd1 vccd1 _10224_/X sky130_fd_sc_hd__buf_4
XANTENNA__09754__A _11222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17820_ _17820_/A vssd1 vssd1 vccd1 vccd1 _19711_/D sky130_fd_sc_hd__clkbuf_1
X_10155_ _09173_/A _10154_/X _10210_/A vssd1 vssd1 vccd1 vccd1 _10155_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12180__A _12180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17751_ _17751_/A _18485_/Q _17751_/C vssd1 vssd1 vccd1 vccd1 _17757_/B sky130_fd_sc_hd__or3_1
X_14963_ _16709_/A vssd1 vssd1 vccd1 vccd1 _16813_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11508__B _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10086_ _10270_/A vssd1 vssd1 vccd1 vccd1 _10167_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10412__B _12482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output137_A _12465_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16702_ _16702_/A vssd1 vssd1 vccd1 vccd1 _16702_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15491__A _15590_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13914_ _13691_/X _13613_/X _13966_/S vssd1 vssd1 vccd1 vccd1 _13914_/X sky130_fd_sc_hd__mux2_1
X_17682_ _17682_/A vssd1 vssd1 vccd1 vccd1 _19673_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14894_ _18473_/Q _18474_/Q _14894_/C vssd1 vssd1 vccd1 vccd1 _14912_/B sky130_fd_sc_hd__and3_1
XFILLER_90_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19421_ _19616_/CLK _19421_/D vssd1 vssd1 vccd1 vccd1 _19421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16633_ _19272_/Q vssd1 vssd1 vccd1 vccd1 _16634_/A sky130_fd_sc_hd__clkbuf_1
X_13845_ _13843_/X _13844_/X _13845_/S vssd1 vssd1 vccd1 vccd1 _13846_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19352_ _19610_/CLK _19352_/D vssd1 vssd1 vccd1 vccd1 _19352_/Q sky130_fd_sc_hd__dfxtp_1
X_16564_ _16564_/A vssd1 vssd1 vccd1 vccd1 _19237_/D sky130_fd_sc_hd__clkbuf_1
X_13776_ _13774_/Y _13775_/X _13776_/S vssd1 vssd1 vccd1 vccd1 _13776_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10988_ _09177_/A _10987_/X _19694_/Q vssd1 vssd1 vccd1 vccd1 _10988_/X sky130_fd_sc_hd__o21a_1
X_18303_ _19788_/CLK _18303_/D vssd1 vssd1 vccd1 vccd1 _18303_/Q sky130_fd_sc_hd__dfxtp_1
X_15515_ _15515_/A vssd1 vssd1 vccd1 vccd1 _18792_/D sky130_fd_sc_hd__clkbuf_1
X_12727_ _12600_/X _12718_/Y _12726_/X _12558_/X _18631_/Q vssd1 vssd1 vccd1 vccd1
+ _12727_/X sky130_fd_sc_hd__a32o_4
X_19283_ _19659_/CLK _19283_/D vssd1 vssd1 vccd1 vccd1 _19283_/Q sky130_fd_sc_hd__dfxtp_1
X_16495_ _16125_/X _19207_/Q _16497_/S vssd1 vssd1 vccd1 vccd1 _16496_/A sky130_fd_sc_hd__mux2_1
X_18234_ _18234_/A vssd1 vssd1 vccd1 vccd1 _18239_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15446_ _18766_/Q _15181_/X _15448_/S vssd1 vssd1 vccd1 vccd1 _15447_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12658_ _12658_/A vssd1 vssd1 vccd1 vccd1 _14648_/A sky130_fd_sc_hd__buf_2
XFILLER_157_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18165_ _18165_/A _18165_/B _18167_/B vssd1 vssd1 vccd1 vccd1 _19842_/D sky130_fd_sc_hd__nor3_1
X_11609_ _11618_/B vssd1 vssd1 vccd1 vccd1 _11940_/A sky130_fd_sc_hd__buf_2
X_15377_ _15377_/A vssd1 vssd1 vccd1 vccd1 _18736_/D sky130_fd_sc_hd__clkbuf_1
X_12589_ _18346_/Q _12643_/A _12674_/A _18400_/Q _12588_/X vssd1 vssd1 vccd1 vccd1
+ _12589_/X sky130_fd_sc_hd__a221o_1
XANTENNA__12355__A _12355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17116_ _17116_/A vssd1 vssd1 vccd1 vccd1 _19457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14328_ _14328_/A _14328_/B vssd1 vssd1 vccd1 vccd1 _14328_/Y sky130_fd_sc_hd__nand2_1
XFILLER_171_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18096_ _18120_/A _18096_/B _18096_/C vssd1 vssd1 vccd1 vccd1 _19818_/D sky130_fd_sc_hd__nor3_1
XFILLER_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17357__S _17363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17047_ _19427_/Q _16718_/X _17047_/S vssd1 vssd1 vccd1 vccd1 _17048_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15666__A _15734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14259_ _18450_/Q _14258_/X _14306_/S vssd1 vssd1 vccd1 vccd1 _14260_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18042__A _18085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12165__A0 _12163_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09664__A _10390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10603__A _10622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ _19549_/CLK _18998_/D vssd1 vssd1 vccd1 vccd1 _18998_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17949_ _19767_/Q _17945_/C _17948_/Y vssd1 vssd1 vccd1 vccd1 _19767_/D sky130_fd_sc_hd__o21a_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19619_ _19833_/CLK _19619_/D vssd1 vssd1 vccd1 vccd1 _19619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10326__S0 _10125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09303_ _09303_/A _09303_/B _09303_/C _09303_/D vssd1 vssd1 vccd1 vccd1 _09624_/B
+ sky130_fd_sc_hd__and4_4
XFILLER_62_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16436__S _16442_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09234_ _19532_/Q _19146_/Q _19596_/Q _18752_/Q _09190_/X _09165_/A vssd1 vssd1 vccd1
+ vccd1 _09235_/B sky130_fd_sc_hd__mux4_1
XFILLER_21_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12928__C1 _12802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09165_ _09165_/A _09165_/B vssd1 vssd1 vccd1 vccd1 _09165_/X sky130_fd_sc_hd__and2_1
XFILLER_148_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09096_ _11337_/A vssd1 vssd1 vccd1 vccd1 _11376_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10954__B2 _18429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17267__S _17269_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11903__A0 _11899_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13096__A _17892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11609__A _11618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09293__B _15134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ _10020_/A _09998_/B vssd1 vssd1 vccd1 vccd1 _09998_/X sky130_fd_sc_hd__or2_1
XFILLER_131_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13105__C1 _13102_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11328__B _11514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11960_ _11847_/X _11958_/X _11959_/X _11560_/X vssd1 vssd1 vccd1 vccd1 _11960_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10911_ _19245_/Q _19016_/Q _18947_/Q _19341_/Q _10909_/X _10910_/X vssd1 vssd1 vccd1
+ vccd1 _10911_/X sky130_fd_sc_hd__mux4_2
XFILLER_56_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11891_ _11886_/X _11890_/Y _11901_/A _11788_/B vssd1 vssd1 vccd1 vccd1 _17870_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13630_ _13630_/A vssd1 vssd1 vccd1 vccd1 _13936_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10842_ _19408_/Q _19184_/Q _19701_/Q _19152_/Q _10648_/S _10785_/X vssd1 vssd1 vccd1
+ vccd1 _10842_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12159__B _13598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09627__A2 _09607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13561_ _13561_/A vssd1 vssd1 vccd1 vccd1 _18424_/D sky130_fd_sc_hd__clkbuf_1
X_10773_ _19249_/Q _19020_/Q _18951_/Q _19345_/Q _10719_/X _10772_/X vssd1 vssd1 vccd1
+ vccd1 _10773_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15300_ _18703_/Q _15184_/X _15300_/S vssd1 vssd1 vccd1 vccd1 _15301_/A sky130_fd_sc_hd__mux2_1
X_12512_ _18417_/Q vssd1 vssd1 vccd1 vccd1 _12766_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10642__B1 _09409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16280_ _16280_/A vssd1 vssd1 vccd1 vccd1 _19112_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13492_ _13492_/A vssd1 vssd1 vccd1 vccd1 _18404_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15231_ _15231_/A vssd1 vssd1 vccd1 vccd1 _18679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12443_ _12505_/A _12345_/X _11941_/Y vssd1 vssd1 vccd1 vccd1 _14332_/B sky130_fd_sc_hd__o21ai_4
XFILLER_60_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15162_ _16664_/A vssd1 vssd1 vccd1 vccd1 _15162_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12374_ _12371_/B _12331_/X _12371_/C _12373_/X _12354_/B vssd1 vssd1 vccd1 vccd1
+ _12374_/X sky130_fd_sc_hd__a311o_1
XFILLER_158_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14113_ _13795_/A _14110_/Y _14112_/X vssd1 vssd1 vccd1 vccd1 _14113_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11325_ _14578_/A _14575_/A _11325_/C _09125_/A vssd1 vssd1 vccd1 vccd1 _11375_/B
+ sky130_fd_sc_hd__or4b_2
XFILLER_4_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16081__S _16081_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15093_ _18623_/Q _15092_/X _15093_/S vssd1 vssd1 vccd1 vccd1 _15094_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12147__B1 _17221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18921_ _19541_/CLK _18921_/D vssd1 vssd1 vccd1 vccd1 _18921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14044_ _13927_/A _14043_/Y _13856_/A vssd1 vssd1 vccd1 vccd1 _14044_/Y sky130_fd_sc_hd__a21oi_1
X_11256_ _11220_/A _11249_/Y _11199_/Y vssd1 vssd1 vccd1 vccd1 _11258_/B sky130_fd_sc_hd__a21oi_2
XFILLER_122_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17086__A0 _16774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10207_ _10210_/A _10204_/X _10206_/X _09988_/A vssd1 vssd1 vccd1 vccd1 _10207_/X
+ sky130_fd_sc_hd__o211a_1
X_11187_ _11187_/A vssd1 vssd1 vccd1 vccd1 _11187_/Y sky130_fd_sc_hd__inv_2
X_18852_ _19534_/CLK _18852_/D vssd1 vssd1 vccd1 vccd1 _18852_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_151_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ _09318_/A _10127_/Y _10133_/X _10137_/Y _09395_/A vssd1 vssd1 vccd1 vccd1
+ _10138_/X sky130_fd_sc_hd__o311a_1
X_17803_ _15165_/X _19704_/Q _17805_/S vssd1 vssd1 vccd1 vccd1 _17804_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13647__A0 _13665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18783_ _19285_/CLK _18783_/D vssd1 vssd1 vccd1 vccd1 _18783_/Q sky130_fd_sc_hd__dfxtp_1
X_15995_ _15995_/A vssd1 vssd1 vccd1 vccd1 _18996_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17734_ _12757_/X _17733_/Y _17734_/S vssd1 vssd1 vccd1 vccd1 _17734_/X sky130_fd_sc_hd__mux2_1
X_10069_ _19617_/Q _19455_/Q _18901_/Q _18671_/Q _10033_/S _09880_/A vssd1 vssd1 vccd1
+ vccd1 _10069_/X sky130_fd_sc_hd__mux4_1
X_14946_ _14958_/A _14946_/B _14946_/C _14946_/D vssd1 vssd1 vccd1 vccd1 _14946_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_36_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17665_ _19670_/Q _17664_/X _17681_/S vssd1 vssd1 vccd1 vccd1 _17666_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14877_ _14877_/A _14877_/B vssd1 vssd1 vccd1 vccd1 _16686_/A sky130_fd_sc_hd__nor2_4
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16616_ _16616_/A vssd1 vssd1 vccd1 vccd1 _19263_/D sky130_fd_sc_hd__clkbuf_1
X_19404_ _19697_/CLK _19404_/D vssd1 vssd1 vccd1 vccd1 _19404_/Q sky130_fd_sc_hd__dfxtp_1
X_13828_ _14173_/A vssd1 vssd1 vccd1 vccd1 _13828_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10881__B1 _12466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17596_ _17596_/A vssd1 vssd1 vccd1 vccd1 _19655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19335_ _19590_/CLK _19335_/D vssd1 vssd1 vccd1 vccd1 _19335_/Q sky130_fd_sc_hd__dfxtp_1
X_16547_ _19230_/Q _15551_/X _16547_/S vssd1 vssd1 vccd1 vccd1 _16548_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13759_ _13757_/X _13758_/X _13759_/S vssd1 vssd1 vccd1 vccd1 _13955_/B sky130_fd_sc_hd__mux2_1
XFILLER_149_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14565__A _14565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19266_ _19589_/CLK _19266_/D vssd1 vssd1 vccd1 vccd1 _19266_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09659__A _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16478_ _16099_/X _19199_/Q _16486_/S vssd1 vssd1 vccd1 vccd1 _16479_/A sky130_fd_sc_hd__mux2_1
X_18217_ _18223_/A _18222_/C vssd1 vssd1 vccd1 vccd1 _18217_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17876__A _17882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15429_ _18758_/Q _15155_/X _15437_/S vssd1 vssd1 vccd1 vccd1 _15430_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19197_ _19647_/CLK _19197_/D vssd1 vssd1 vccd1 vccd1 _19197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_76_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18148_ _19836_/Q _19835_/Q _18148_/C vssd1 vssd1 vccd1 vccd1 _18150_/B sky130_fd_sc_hd__and3_1
XFILLER_163_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18079_ _18079_/A vssd1 vssd1 vccd1 vccd1 _18086_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09921_ _09905_/A _09920_/X _09231_/X vssd1 vssd1 vccd1 vccd1 _09921_/X sky130_fd_sc_hd__o21a_1
XFILLER_104_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09394__A _09394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11036__S1 _10960_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09852_ _09992_/A _09852_/B vssd1 vssd1 vccd1 vccd1 _09852_/X sky130_fd_sc_hd__or2_1
XFILLER_112_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11148__B _12497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09783_ _09783_/A vssd1 vssd1 vccd1 vccd1 _09783_/X sky130_fd_sc_hd__buf_2
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15335__S _15337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13363__B _13363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10321__C1 _09562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16955__A _16977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16166__S _16172_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09217_ _09217_/A vssd1 vssd1 vccd1 vccd1 _09217_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__16690__A _16722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09148_ _09841_/A vssd1 vssd1 vccd1 vccd1 _09149_/A sky130_fd_sc_hd__buf_4
XFILLER_147_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09079_ _18568_/Q vssd1 vssd1 vccd1 vccd1 _09125_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11110_ _18862_/Q _19320_/Q _11110_/S vssd1 vssd1 vccd1 vccd1 _11110_/X sky130_fd_sc_hd__mux2_1
X_12090_ _19744_/Q vssd1 vssd1 vccd1 vccd1 _12095_/A sky130_fd_sc_hd__buf_4
XFILLER_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11041_ _11041_/A _11041_/B vssd1 vssd1 vccd1 vccd1 _11041_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10243__A _10451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10786__S0 _10711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14800_ _14795_/Y _14827_/C _14798_/X _14980_/A vssd1 vssd1 vccd1 vccd1 _14800_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _14940_/X _18900_/Q _15780_/S vssd1 vssd1 vccd1 vccd1 _15781_/A sky130_fd_sc_hd__mux2_1
X_12992_ _12993_/A _12993_/C _18311_/Q vssd1 vssd1 vccd1 vccd1 _12994_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__11104__A1 _09434_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12301__B1 _19752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14731_ _14731_/A vssd1 vssd1 vccd1 vccd1 _18587_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input13_A io_dbus_rdata[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10389__S _10389_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11943_ _11470_/A _11941_/Y _11942_/Y vssd1 vssd1 vccd1 vccd1 _11943_/X sky130_fd_sc_hd__o21a_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _17450_/A vssd1 vssd1 vccd1 vccd1 _19590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14662_ _14662_/A vssd1 vssd1 vccd1 vccd1 _18573_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ _11745_/A _11783_/B _11811_/Y vssd1 vssd1 vccd1 vccd1 _11874_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16401_ _16401_/A vssd1 vssd1 vccd1 vccd1 _19165_/D sky130_fd_sc_hd__clkbuf_1
X_13613_ _13602_/X _13611_/X _13759_/S vssd1 vssd1 vccd1 vccd1 _13613_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10825_ _10866_/A _10825_/B vssd1 vssd1 vccd1 vccd1 _10825_/X sky130_fd_sc_hd__or2_1
X_17381_ _16832_/X _19560_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _17382_/A sky130_fd_sc_hd__mux2_1
X_14593_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14593_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19120_ _19614_/CLK _19120_/D vssd1 vssd1 vccd1 vccd1 _19120_/Q sky130_fd_sc_hd__dfxtp_1
X_16332_ _16099_/X _19135_/Q _16340_/S vssd1 vssd1 vccd1 vccd1 _16333_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13544_ _13563_/A vssd1 vssd1 vccd1 vccd1 _13560_/A sky130_fd_sc_hd__clkbuf_1
X_10756_ _10750_/A _10753_/X _10755_/X _09225_/A vssd1 vssd1 vccd1 vccd1 _10756_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12617__B _12617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10091__A1 _10107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19051_ _19614_/CLK _19051_/D vssd1 vssd1 vccd1 vccd1 _19051_/Q sky130_fd_sc_hd__dfxtp_1
X_16263_ _16263_/A vssd1 vssd1 vccd1 vccd1 _19104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13475_ _18397_/Q _13294_/X _13475_/S vssd1 vssd1 vccd1 vccd1 _13476_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10687_ _10752_/A _10687_/B vssd1 vssd1 vccd1 vccd1 _10687_/X sky130_fd_sc_hd__or2_1
XANTENNA__10630__A3 _10629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16804__S _16807_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18002_ _19785_/Q _18000_/B _18001_/Y vssd1 vssd1 vccd1 vccd1 _19785_/D sky130_fd_sc_hd__o21a_1
X_15214_ _18674_/Q _15213_/X _15217_/S vssd1 vssd1 vccd1 vccd1 _15215_/A sky130_fd_sc_hd__mux2_1
X_12426_ _12426_/A _14324_/B vssd1 vssd1 vccd1 vccd1 _12426_/X sky130_fd_sc_hd__or2_1
X_16194_ _16112_/X _19070_/Q _16194_/S vssd1 vssd1 vccd1 vccd1 _16195_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14109__A1 _14126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15145_ _15145_/A vssd1 vssd1 vccd1 vccd1 _18652_/D sky130_fd_sc_hd__clkbuf_1
X_12357_ _12371_/C _12357_/B vssd1 vssd1 vccd1 vccd1 _14284_/A sky130_fd_sc_hd__xnor2_4
XFILLER_154_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11308_ _13568_/A _13568_/B _11287_/X vssd1 vssd1 vccd1 vccd1 _11736_/A sky130_fd_sc_hd__or3b_2
X_15076_ _16844_/A vssd1 vssd1 vccd1 vccd1 _15076_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12288_ _12262_/A _14241_/B _12287_/X vssd1 vssd1 vccd1 vccd1 _12288_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_141_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12352__B _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18904_ _19395_/CLK _18904_/D vssd1 vssd1 vccd1 vccd1 _18904_/Q sky130_fd_sc_hd__dfxtp_1
X_14027_ _13942_/A _14024_/Y _14026_/Y _13711_/B vssd1 vssd1 vccd1 vccd1 _14027_/X
+ sky130_fd_sc_hd__a211o_1
X_11239_ _11239_/A vssd1 vssd1 vccd1 vccd1 _11239_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10777__S0 _10934_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18835_ _19715_/CLK _18835_/D vssd1 vssd1 vccd1 vccd1 _18835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15978_ _15978_/A vssd1 vssd1 vccd1 vccd1 _18988_/D sky130_fd_sc_hd__clkbuf_1
X_18766_ _19610_/CLK _18766_/D vssd1 vssd1 vccd1 vccd1 _18766_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09839__A2 _09817_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17717_ _12656_/B _17716_/Y _17734_/S vssd1 vssd1 vccd1 vccd1 _17717_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14929_ _16803_/A vssd1 vssd1 vccd1 vccd1 _14929_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18697_ _19638_/CLK _18697_/D vssd1 vssd1 vccd1 vccd1 _18697_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10600__B _12474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17370__S _17374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17648_ _17648_/A vssd1 vssd1 vccd1 vccd1 _19667_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17579_ _19648_/Q _16806_/A _17579_/S vssd1 vssd1 vccd1 vccd1 _17580_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19318_ _19608_/CLK _19318_/D vssd1 vssd1 vccd1 vccd1 _19318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19249_ _19703_/CLK _19249_/D vssd1 vssd1 vccd1 vccd1 _19249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18214__B _18214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09870__S1 _09869_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12262__B _12262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09904_ _19652_/Q _19069_/Q _19106_/Q _18712_/Q _09782_/X _09763_/X vssd1 vssd1 vccd1
+ vccd1 _09905_/B sky130_fd_sc_hd__mux4_2
XFILLER_120_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09835_ _09879_/A _09834_/X _09320_/A vssd1 vssd1 vccd1 vccd1 _09835_/X sky130_fd_sc_hd__o21a_1
XFILLER_112_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input5_A io_dbus_rdata[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09766_ _18873_/Q _19331_/Q _10010_/S vssd1 vssd1 vccd1 vccd1 _09767_/B sky130_fd_sc_hd__mux2_1
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13087__B2 _18626_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14189__B _14192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ _09697_/A vssd1 vssd1 vccd1 vccd1 _10103_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__17222__A0 _18450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17280__S _17280_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10610_ _10830_/A vssd1 vssd1 vccd1 vccd1 _10750_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11590_ _11618_/A vssd1 vssd1 vccd1 vccd1 _13625_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15536__A0 _18799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14339__A1 _18457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10541_ _18859_/Q _19317_/Q _10604_/S vssd1 vssd1 vccd1 vccd1 _10541_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10238__A _10238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13260_ _13438_/B vssd1 vssd1 vccd1 vccd1 _13295_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10472_ _11099_/A _10469_/X _10471_/X _09227_/A vssd1 vssd1 vccd1 vccd1 _10472_/X
+ sky130_fd_sc_hd__o211a_1
X_12211_ _12185_/A _12185_/B _12182_/A vssd1 vssd1 vccd1 vccd1 _12212_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__13562__A2 _13536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13191_ _19474_/Q _12741_/X _13189_/X _13190_/X vssd1 vssd1 vccd1 vccd1 _13191_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12453__A _19690_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ _12142_/A vssd1 vssd1 vccd1 vccd1 _12142_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17455__S _17457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12073_ _11980_/A _12070_/X _12071_/X _12072_/X vssd1 vssd1 vccd1 vccd1 _12073_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16950_ _16950_/A vssd1 vssd1 vccd1 vccd1 _19383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10759__S0 _10836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15901_ _15901_/A vssd1 vssd1 vccd1 vccd1 _18953_/D sky130_fd_sc_hd__clkbuf_1
X_11024_ _11619_/A _12460_/A vssd1 vssd1 vccd1 vccd1 _11024_/X sky130_fd_sc_hd__or2_1
XFILLER_77_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16881_ _16881_/A vssd1 vssd1 vccd1 vccd1 _19353_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11876__A2 _13658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_24_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15832_ _15878_/S vssd1 vssd1 vccd1 vccd1 _15841_/S sky130_fd_sc_hd__buf_2
X_18620_ _18623_/CLK _18620_/D vssd1 vssd1 vccd1 vccd1 _18620_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_77_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11089__B1 _09454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ _19732_/CLK _18551_/D vssd1 vssd1 vccd1 vccd1 _18551_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15763_ _14847_/X _18892_/Q _15769_/S vssd1 vssd1 vccd1 vccd1 _15764_/A sky130_fd_sc_hd__mux2_1
X_12975_ _12984_/D vssd1 vssd1 vccd1 vccd1 _12982_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11184__S0 _10129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14714_ _16743_/A vssd1 vssd1 vccd1 vccd1 _14714_/X sky130_fd_sc_hd__buf_2
X_17502_ _17502_/A vssd1 vssd1 vccd1 vccd1 _19613_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18482_ _18482_/CLK _18482_/D vssd1 vssd1 vccd1 vccd1 _18482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11926_ _11930_/B vssd1 vssd1 vccd1 vccd1 _11926_/Y sky130_fd_sc_hd__clkinv_2
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15694_ _15694_/A vssd1 vssd1 vccd1 vccd1 _18861_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09701__S _09701_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _16803_/X _19583_/Q _17435_/S vssd1 vssd1 vccd1 vccd1 _17434_/A sky130_fd_sc_hd__mux2_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _14672_/A _14645_/B vssd1 vssd1 vccd1 vccd1 _18568_/D sky130_fd_sc_hd__nor2_1
X_11857_ _11758_/X _11888_/D _13215_/A vssd1 vssd1 vccd1 vccd1 _11857_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12628__A _12628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17364_ _17364_/A vssd1 vssd1 vccd1 vccd1 _19552_/D sky130_fd_sc_hd__clkbuf_1
X_10808_ _10803_/A _10804_/X _10807_/X _10728_/X vssd1 vssd1 vccd1 vccd1 _10808_/X
+ sky130_fd_sc_hd__o211a_1
X_14576_ _18547_/Q _14564_/X _14575_/X _14573_/X vssd1 vssd1 vccd1 vccd1 _18547_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17516__A1 _16715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11788_ _19733_/Q _11788_/B vssd1 vssd1 vccd1 vccd1 _11803_/A sky130_fd_sc_hd__or2_1
XFILLER_159_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19103_ _19810_/CLK _19103_/D vssd1 vssd1 vccd1 vccd1 _19103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16315_ _16315_/A vssd1 vssd1 vccd1 vccd1 _19127_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13527_ _11470_/A _13527_/B _13527_/C vssd1 vssd1 vccd1 vccd1 _13527_/X sky130_fd_sc_hd__and3b_1
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17295_ _17295_/A vssd1 vssd1 vccd1 vccd1 _19521_/D sky130_fd_sc_hd__clkbuf_1
X_10739_ _10739_/A vssd1 vssd1 vccd1 vccd1 _10740_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_174_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10148__A _18445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19034_ _19810_/CLK _19034_/D vssd1 vssd1 vccd1 vccd1 _19034_/Q sky130_fd_sc_hd__dfxtp_1
X_16246_ _16080_/X _19097_/Q _16246_/S vssd1 vssd1 vccd1 vccd1 _16247_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ _18389_/Q _13212_/X _13464_/S vssd1 vssd1 vccd1 vccd1 _13459_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12409_ _19757_/Q _12410_/B vssd1 vssd1 vccd1 vccd1 _12434_/B sky130_fd_sc_hd__and2_1
XFILLER_126_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16177_ _16087_/X _19062_/Q _16183_/S vssd1 vssd1 vccd1 vccd1 _16178_/A sky130_fd_sc_hd__mux2_1
X_13389_ _13354_/X _13387_/X _13388_/X _13350_/X vssd1 vssd1 vccd1 vccd1 _18377_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput105 _09106_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_ld_type[0] sky130_fd_sc_hd__buf_2
XFILLER_142_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput116 _12482_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[14] sky130_fd_sc_hd__buf_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput127 _12497_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[24] sky130_fd_sc_hd__buf_2
Xoutput138 _12467_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[5] sky130_fd_sc_hd__buf_2
X_15128_ _18646_/Q _15123_/X _15125_/X _09688_/A vssd1 vssd1 vccd1 vccd1 _18646_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput149 _17882_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[14] sky130_fd_sc_hd__buf_2
XFILLER_114_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14502__A1 _19759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15059_ _18488_/Q _15059_/B vssd1 vssd1 vccd1 vccd1 _15059_/X sky130_fd_sc_hd__or2_1
XFILLER_99_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09672__A _10401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19867_ _19871_/CLK _19867_/D vssd1 vssd1 vccd1 vccd1 _19867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11707__A _19731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ _19626_/Q _19464_/Q _18910_/Q _18680_/Q _09344_/A _11189_/A vssd1 vssd1 vccd1
+ vccd1 _09620_/X sky130_fd_sc_hd__mux4_2
X_18818_ _18818_/CLK _18818_/D vssd1 vssd1 vccd1 vccd1 _18818_/Q sky130_fd_sc_hd__dfxtp_1
X_19798_ _19798_/CLK _19798_/D vssd1 vssd1 vccd1 vccd1 _19798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09551_ _10432_/A vssd1 vssd1 vccd1 vccd1 _10309_/A sky130_fd_sc_hd__buf_2
X_18749_ _19271_/CLK _18749_/D vssd1 vssd1 vccd1 vccd1 _18749_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11175__S0 _10129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09482_ _09482_/A vssd1 vssd1 vccd1 vccd1 _09662_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17755__A1 _19686_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18225__A _18225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18180__A1 _19847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09582__A _11110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09818_ _19267_/Q _19038_/Q _18969_/Q _19363_/Q _09803_/X _09875_/A vssd1 vssd1 vccd1
+ vccd1 _09819_/B sky130_fd_sc_hd__mux4_1
XFILLER_74_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09749_ _10127_/A _09748_/X _09621_/X vssd1 vssd1 vccd1 vccd1 _09749_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_28_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14928__A _16699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17304__A _17304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _14431_/A vssd1 vssd1 vccd1 vccd1 _14516_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__13480__A1 _12559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17746__A1 _19684_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10913__S0 _10909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _19662_/Q _12390_/B vssd1 vssd1 vccd1 vccd1 _11711_/X sky130_fd_sc_hd__or2_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12691_ _13536_/A vssd1 vssd1 vccd1 vccd1 _14577_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14430_ _14430_/A vssd1 vssd1 vccd1 vccd1 _18489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _13526_/A _13583_/A _11642_/C vssd1 vssd1 vccd1 vccd1 _13571_/B sky130_fd_sc_hd__or3_1
XFILLER_168_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14361_ _18465_/Q _18497_/Q _14367_/S vssd1 vssd1 vccd1 vccd1 _14362_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11573_ _11325_/C _11337_/A _11484_/A _11484_/B _11472_/A vssd1 vssd1 vccd1 vccd1
+ _11735_/S sky130_fd_sc_hd__o2111a_1
XFILLER_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16100_ _16116_/A vssd1 vssd1 vccd1 vccd1 _16113_/S sky130_fd_sc_hd__buf_4
XANTENNA__10141__S1 _10186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput18 io_dbus_rdata[25] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_2
X_13312_ _13312_/A _13319_/B vssd1 vssd1 vccd1 vccd1 _13312_/X sky130_fd_sc_hd__or2_1
XFILLER_156_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17080_ _16765_/X _19441_/Q _17086_/S vssd1 vssd1 vccd1 vccd1 _17081_/A sky130_fd_sc_hd__mux2_1
Xinput29 io_dbus_rdata[6] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_4
X_10524_ _10524_/A _10524_/B vssd1 vssd1 vccd1 vccd1 _10524_/X sky130_fd_sc_hd__or2_1
XANTENNA__09757__A _10257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14292_ _14150_/X _13918_/X _14291_/X _13823_/X vssd1 vssd1 vccd1 vccd1 _14292_/X
+ sky130_fd_sc_hd__a211o_1
X_16031_ _15076_/X _19013_/Q _16031_/S vssd1 vssd1 vccd1 vccd1 _16032_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09739__A1 _11178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13243_ _19769_/Q _12753_/X _13242_/X vssd1 vssd1 vccd1 vccd1 _14813_/D sky130_fd_sc_hd__a21o_1
XFILLER_6_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10455_ _10395_/A _10454_/X _09314_/A vssd1 vssd1 vccd1 vccd1 _10455_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09834__S1 _09810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ _19663_/Q _13251_/A _13154_/B _18387_/Q vssd1 vssd1 vccd1 vccd1 _13174_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10386_ _10400_/A _10386_/B vssd1 vssd1 vccd1 vccd1 _10386_/Y sky130_fd_sc_hd__nor2_1
X_12125_ _19745_/Q _12116_/X _12121_/Y _12124_/Y vssd1 vssd1 vccd1 vccd1 _17888_/B
+ sky130_fd_sc_hd__o22a_1
X_17982_ _17991_/A _17988_/C vssd1 vssd1 vccd1 vccd1 _17982_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14496__A0 _18518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13299__B2 _19839_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19721_ _19721_/CLK _19721_/D vssd1 vssd1 vccd1 vccd1 _19721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16933_ _16990_/S vssd1 vssd1 vccd1 vccd1 _16942_/S sky130_fd_sc_hd__buf_2
X_12056_ _12131_/C vssd1 vssd1 vccd1 vccd1 _14140_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_104_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _11003_/X _11005_/X _11006_/X _11060_/A _10774_/A vssd1 vssd1 vccd1 vccd1
+ _11012_/B sky130_fd_sc_hd__o221a_1
XFILLER_77_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19652_ _19718_/CLK _19652_/D vssd1 vssd1 vccd1 vccd1 _19652_/Q sky130_fd_sc_hd__dfxtp_1
X_16864_ _16864_/A vssd1 vssd1 vccd1 vccd1 _19345_/D sky130_fd_sc_hd__clkbuf_1
X_18603_ _19645_/CLK _18603_/D vssd1 vssd1 vccd1 vccd1 _18603_/Q sky130_fd_sc_hd__dfxtp_1
X_15815_ _14740_/X _18915_/Q _15819_/S vssd1 vssd1 vccd1 vccd1 _15816_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16795_ _16793_/X _19322_/Q _16807_/S vssd1 vssd1 vccd1 vccd1 _16796_/A sky130_fd_sc_hd__mux2_1
X_19583_ _19714_/CLK _19583_/D vssd1 vssd1 vccd1 vccd1 _19583_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10150__B _12488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18534_ _18567_/CLK _18534_/D vssd1 vssd1 vccd1 vccd1 _18534_/Q sky130_fd_sc_hd__dfxtp_1
X_15746_ _15746_/A vssd1 vssd1 vccd1 vccd1 _18884_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12958_ _12983_/A _12958_/B _12959_/B vssd1 vssd1 vccd1 vccd1 _18296_/D sky130_fd_sc_hd__nor3_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13471__A1 _12727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10285__A1 _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11909_ _11885_/X _11907_/X _11936_/B _11625_/A vssd1 vssd1 vccd1 vccd1 _11909_/X
+ sky130_fd_sc_hd__a31o_1
X_15677_ _15734_/S vssd1 vssd1 vccd1 vccd1 _15686_/S sky130_fd_sc_hd__buf_2
X_18465_ _19693_/CLK _18465_/D vssd1 vssd1 vccd1 vccd1 _18465_/Q sky130_fd_sc_hd__dfxtp_1
X_12889_ _18276_/Q vssd1 vssd1 vccd1 vccd1 _12895_/C sky130_fd_sc_hd__clkbuf_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12358__A _14284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10380__S1 _09554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14628_ _14654_/A _14628_/B vssd1 vssd1 vccd1 vccd1 _14629_/A sky130_fd_sc_hd__and2_1
X_17416_ _16777_/X _19575_/Q _17424_/S vssd1 vssd1 vccd1 vccd1 _17417_/A sky130_fd_sc_hd__mux2_1
X_18396_ _19687_/CLK _18396_/D vssd1 vssd1 vccd1 vccd1 _18396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17347_ _17347_/A vssd1 vssd1 vccd1 vccd1 _19544_/D sky130_fd_sc_hd__clkbuf_1
X_14559_ _14559_/A _14559_/B vssd1 vssd1 vccd1 vccd1 _14559_/X sky130_fd_sc_hd__or2_1
XFILLER_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13774__A2 _13720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16264__S _16268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18045__A _18077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17278_ _19514_/Q _16683_/X _17280_/S vssd1 vssd1 vccd1 vccd1 _17279_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19017_ _19568_/CLK _19017_/D vssd1 vssd1 vccd1 vccd1 _19017_/Q sky130_fd_sc_hd__dfxtp_1
X_16229_ _16055_/X _19089_/Q _16235_/S vssd1 vssd1 vccd1 vccd1 _16230_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15920__A0 _14918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17884__A _17890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17095__S _17097_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17823__S _17827_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10341__A _11185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09603_ _09603_/A vssd1 vssd1 vccd1 vccd1 _09610_/A sky130_fd_sc_hd__buf_2
XFILLER_83_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15343__S _15351_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09534_ _11202_/A _12504_/A vssd1 vssd1 vccd1 vccd1 _11203_/A sky130_fd_sc_hd__and2_2
XANTENNA__13462__A1 _13230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15739__A0 _14714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09465_ _11097_/A _09465_/B vssd1 vssd1 vccd1 vccd1 _09465_/X sky130_fd_sc_hd__or2_1
XFILLER_145_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09396_ _09320_/X _09366_/Y _09371_/X _09388_/Y _09395_/X vssd1 vssd1 vccd1 vccd1
+ _09396_/X sky130_fd_sc_hd__o311a_1
XANTENNA__10028__B2 _18447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18153__A1 _19838_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12715__B _12715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13099__A input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16902__S _16902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10240_ _18866_/Q _19324_/Q _10401_/A vssd1 vssd1 vccd1 vccd1 _10241_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17664__A0 _12713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16467__A1 _19194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10171_ _09278_/A _10161_/X _10170_/X _09285_/A _18444_/Q vssd1 vssd1 vccd1 vccd1
+ _10196_/A sky130_fd_sc_hd__a32o_4
XFILLER_121_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12731__A _12731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13930_ _13926_/X _13930_/B vssd1 vssd1 vccd1 vccd1 _13931_/C sky130_fd_sc_hd__and2b_1
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13861_ _13745_/X _13665_/X _14323_/A vssd1 vssd1 vccd1 vccd1 _13862_/C sky130_fd_sc_hd__a21oi_1
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16349__S _16351_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14658__A _14677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15600_ _15600_/A vssd1 vssd1 vccd1 vccd1 _18819_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12812_ _18225_/A vssd1 vssd1 vccd1 vccd1 _12844_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16580_ _16580_/A vssd1 vssd1 vccd1 vccd1 _19245_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13453__A1 _13182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13792_ _13888_/S vssd1 vssd1 vccd1 vccd1 _13839_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_16_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15531_ _15531_/A vssd1 vssd1 vccd1 vccd1 _18797_/D sky130_fd_sc_hd__clkbuf_1
X_12743_ _13154_/B vssd1 vssd1 vccd1 vccd1 _12743_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18250_ _18250_/A _18250_/B vssd1 vssd1 vccd1 vccd1 _18250_/Y sky130_fd_sc_hd__nor2_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15462_ _18773_/Q _15203_/X _15470_/S vssd1 vssd1 vccd1 vccd1 _15463_/A sky130_fd_sc_hd__mux2_1
X_12674_ _12674_/A vssd1 vssd1 vccd1 vccd1 _13428_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _18444_/Q _12617_/B _17201_/S vssd1 vssd1 vccd1 vccd1 _17201_/X sky130_fd_sc_hd__mux2_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _18483_/Q _18515_/Q _14424_/S vssd1 vssd1 vccd1 vccd1 _14414_/A sky130_fd_sc_hd__mux2_1
X_18181_ _19847_/Q _18183_/C _18180_/Y vssd1 vssd1 vccd1 vccd1 _19847_/D sky130_fd_sc_hd__o21a_1
X_11625_ _11625_/A vssd1 vssd1 vccd1 vccd1 _11997_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15489__A _16503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15393_ _18744_/Q _15213_/X _15395_/S vssd1 vssd1 vccd1 vccd1 _15394_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18144__A1 _19834_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17132_ _16841_/X _19465_/Q _17134_/S vssd1 vssd1 vccd1 vccd1 _17133_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14824__C _14824_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09487__A _18977_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14344_ _14344_/A vssd1 vssd1 vccd1 vccd1 _18459_/D sky130_fd_sc_hd__clkbuf_1
X_11556_ _11556_/A vssd1 vssd1 vccd1 vccd1 _12469_/B sky130_fd_sc_hd__buf_2
XFILLER_156_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10507_ _11082_/B _12478_/B vssd1 vssd1 vccd1 vccd1 _11242_/B sky130_fd_sc_hd__or2b_1
XANTENNA__14705__A1 _13134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17063_ _17063_/A vssd1 vssd1 vccd1 vccd1 _19434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14275_ _13796_/A _14276_/B _14273_/X _14274_/X vssd1 vssd1 vccd1 vccd1 _14275_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_11487_ _13977_/A vssd1 vssd1 vccd1 vccd1 _14250_/A sky130_fd_sc_hd__clkbuf_2
X_16014_ _14986_/X _19005_/Q _16016_/S vssd1 vssd1 vccd1 vccd1 _16015_/A sky130_fd_sc_hd__mux2_1
X_13226_ _19864_/Q _12604_/X _12584_/X _18140_/B _13225_/X vssd1 vssd1 vccd1 vccd1
+ _13226_/X sky130_fd_sc_hd__a221o_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14181__A2 _14176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10438_ _10438_/A _10438_/B vssd1 vssd1 vccd1 vccd1 _10438_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13157_ _12734_/A _13166_/A _15242_/B _12641_/A vssd1 vssd1 vccd1 vccd1 _13157_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_98_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _19417_/Q _19193_/Q _19710_/Q _19161_/Q _09632_/A _10368_/X vssd1 vssd1 vccd1
+ vccd1 _10369_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12108_ _14168_/A _12108_/B vssd1 vssd1 vccd1 vccd1 _12111_/A sky130_fd_sc_hd__xnor2_1
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15130__A1 hold3/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17965_ _19773_/Q _17965_/B vssd1 vssd1 vccd1 vccd1 _17971_/C sky130_fd_sc_hd__and2_1
X_13088_ _13088_/A vssd1 vssd1 vccd1 vccd1 _13110_/A sky130_fd_sc_hd__clkbuf_4
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15130__B2 _11200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13141__B1 _13154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17407__A0 _16765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19704_ _19704_/CLK _19704_/D vssd1 vssd1 vccd1 vccd1 _19704_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15952__A _18207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12039_ _11978_/A _11978_/B _12013_/A _12038_/X vssd1 vssd1 vccd1 vccd1 _12040_/B
+ sky130_fd_sc_hd__a31o_2
X_16916_ _16916_/A vssd1 vssd1 vccd1 vccd1 _19369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17896_ _19748_/Q _17886_/X _12194_/X _12200_/X _17895_/X vssd1 vssd1 vccd1 vccd1
+ _19748_/D sky130_fd_sc_hd__o221a_1
XFILLER_65_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19635_ _19635_/CLK _19635_/D vssd1 vssd1 vccd1 vccd1 _19635_/Q sky130_fd_sc_hd__dfxtp_1
X_16847_ _16847_/A _16847_/B vssd1 vssd1 vccd1 vccd1 _16904_/A sky130_fd_sc_hd__nor2_4
XFILLER_168_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14568__A _14568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11691__S _15095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19566_ _19697_/CLK _19566_/D vssd1 vssd1 vccd1 vccd1 _19566_/Q sky130_fd_sc_hd__dfxtp_1
X_16778_ _16845_/S vssd1 vssd1 vccd1 vccd1 _16791_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__14287__B _14289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10258__A1 _09173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18517_ _18548_/CLK _18517_/D vssd1 vssd1 vccd1 vccd1 _18517_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15729_ _15729_/A vssd1 vssd1 vccd1 vccd1 _18877_/D sky130_fd_sc_hd__clkbuf_1
X_19497_ _19786_/CLK _19497_/D vssd1 vssd1 vccd1 vccd1 _19497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09250_ _09217_/X _09235_/X _09237_/X _09241_/X _09249_/X vssd1 vssd1 vccd1 vccd1
+ _09250_/X sky130_fd_sc_hd__a311o_1
X_18448_ _18632_/CLK _18448_/D vssd1 vssd1 vccd1 vccd1 _18448_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_166_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09181_ _09549_/A vssd1 vssd1 vccd1 vccd1 _11099_/A sky130_fd_sc_hd__clkbuf_4
X_18379_ _19690_/CLK _18379_/D vssd1 vssd1 vccd1 vccd1 _18379_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_146_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17646__A0 _13230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10770__S _10770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15121__B2 _10003_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11694__A0 _12463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14478__A _14591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10249__A1 _11119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09517_ _09517_/A vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__buf_2
XFILLER_25_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16693__A _16693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10010__S _10010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _18616_/Q _19305_/Q _09448_/S vssd1 vssd1 vccd1 vccd1 _09448_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14935__A1 _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09379_ _10395_/A vssd1 vssd1 vccd1 vccd1 _10226_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_138_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12726__A _18631_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11410_ _18544_/Q vssd1 vssd1 vccd1 vccd1 _12533_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__11630__A _12715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15102__A _15116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12390_ _19687_/Q _12390_/B vssd1 vssd1 vccd1 vccd1 _12390_/X sky130_fd_sc_hd__or2_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12445__B _12446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11341_ _11344_/A _11375_/B vssd1 vssd1 vccd1 vccd1 _11372_/A sky130_fd_sc_hd__nor2_2
XFILLER_125_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14060_ _13714_/X _14062_/B _14058_/X _14059_/X vssd1 vssd1 vccd1 vccd1 _14060_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15360__A1 _15165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11272_ _11272_/A vssd1 vssd1 vccd1 vccd1 _11272_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12174__A1 _12489_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ _17993_/A vssd1 vssd1 vccd1 vccd1 _13011_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17637__A0 _19665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10223_ _10581_/S vssd1 vssd1 vccd1 vccd1 _10486_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09754__B _12500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12461__A _12461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input43_A io_ibus_inst[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15112__A1 _18634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ _18867_/Q _19325_/Q _10154_/S vssd1 vssd1 vccd1 vccd1 _10154_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15112__B2 _11135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17750_ _17750_/A vssd1 vssd1 vccd1 vccd1 _19685_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14962_ _14811_/X _14957_/Y _14959_/X _14961_/X vssd1 vssd1 vccd1 vccd1 _16709_/A
+ sky130_fd_sc_hd__o31a_4
XFILLER_59_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10085_ _10262_/A vssd1 vssd1 vccd1 vccd1 _10270_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09770__A _09783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16701_ _16701_/A vssd1 vssd1 vccd1 vccd1 _19293_/D sky130_fd_sc_hd__clkbuf_1
X_13913_ _13684_/X _13664_/X _13913_/S vssd1 vssd1 vccd1 vccd1 _13913_/X sky130_fd_sc_hd__mux2_1
X_17681_ _19673_/Q _17680_/X _17681_/S vssd1 vssd1 vccd1 vccd1 _17682_/A sky130_fd_sc_hd__mux2_1
X_14893_ _14893_/A vssd1 vssd1 vccd1 vccd1 _14969_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19420_ _19635_/CLK _19420_/D vssd1 vssd1 vccd1 vccd1 _19420_/Q sky130_fd_sc_hd__dfxtp_1
X_16632_ _16632_/A vssd1 vssd1 vccd1 vccd1 _19271_/D sky130_fd_sc_hd__clkbuf_1
X_13844_ _13602_/X _13626_/X _13879_/S vssd1 vssd1 vccd1 vccd1 _13844_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12229__A2 _14216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19351_ _19710_/CLK _19351_/D vssd1 vssd1 vccd1 vccd1 _19351_/Q sky130_fd_sc_hd__dfxtp_1
X_16563_ _19237_/Q _15574_/X _16569_/S vssd1 vssd1 vccd1 vccd1 _16564_/A sky130_fd_sc_hd__mux2_1
X_13775_ _13647_/X _13642_/X _13775_/S vssd1 vssd1 vccd1 vccd1 _13775_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16807__S _16807_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10987_ _19404_/Q _19180_/Q _19697_/Q _19148_/Q _10905_/S _10739_/A vssd1 vssd1 vccd1
+ vccd1 _10987_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18302_ _19856_/CLK _18302_/D vssd1 vssd1 vccd1 vccd1 _18302_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15711__S _15719_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12726_ _18631_/Q _12726_/B vssd1 vssd1 vccd1 vccd1 _12726_/X sky130_fd_sc_hd__or2_1
X_15514_ _18792_/Q _15513_/X _15520_/S vssd1 vssd1 vccd1 vccd1 _15515_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19282_ _19537_/CLK _19282_/D vssd1 vssd1 vccd1 vccd1 _19282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16494_ _16494_/A vssd1 vssd1 vccd1 vccd1 _19206_/D sky130_fd_sc_hd__clkbuf_1
X_18233_ _19865_/Q _18230_/A _18232_/Y vssd1 vssd1 vccd1 vccd1 _19865_/D sky130_fd_sc_hd__o21a_1
XFILLER_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15445_ _15445_/A vssd1 vssd1 vccd1 vccd1 _18765_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14926__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12657_ _18336_/Q _12574_/X _12575_/X _12656_/X vssd1 vssd1 vccd1 vccd1 _18336_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11608_ _11686_/A _11686_/B _13587_/B _11686_/D vssd1 vssd1 vccd1 vccd1 _11618_/B
+ sky130_fd_sc_hd__and4_2
X_18164_ _19842_/Q _19841_/Q _18164_/C vssd1 vssd1 vccd1 vccd1 _18167_/B sky130_fd_sc_hd__and3_1
X_15376_ _18736_/Q _15187_/X _15384_/S vssd1 vssd1 vccd1 vccd1 _15377_/A sky130_fd_sc_hd__mux2_1
X_12588_ _19676_/Q _12539_/A _13222_/S _19486_/Q vssd1 vssd1 vccd1 vccd1 _12588_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17115_ _16816_/X _19457_/Q _17119_/S vssd1 vssd1 vccd1 vccd1 _17116_/A sky130_fd_sc_hd__mux2_1
X_14327_ _14150_/X _13782_/X _14326_/X _13823_/X vssd1 vssd1 vccd1 vccd1 _14327_/X
+ sky130_fd_sc_hd__a211o_1
X_18095_ _18094_/A _18094_/C _19818_/Q vssd1 vssd1 vccd1 vccd1 _18096_/C sky130_fd_sc_hd__a21oi_1
X_11539_ _14173_/A _11539_/B _11538_/X vssd1 vssd1 vccd1 vccd1 _11539_/X sky130_fd_sc_hd__or3b_1
XFILLER_172_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17046_ _17046_/A vssd1 vssd1 vccd1 vccd1 _19426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14258_ _12290_/X _14102_/X _14257_/X vssd1 vssd1 vccd1 vccd1 _14258_/X sky130_fd_sc_hd__a21bo_1
XFILLER_172_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17628__A0 _13197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13209_ _19830_/Q _12736_/A _13207_/X _13208_/X vssd1 vssd1 vccd1 vccd1 _13209_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_174_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _14332_/A _14192_/A vssd1 vssd1 vccd1 vccd1 _14189_/X sky130_fd_sc_hd__or2_1
XFILLER_152_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11912__A1 _12476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15103__A1 _18628_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10271__S0 _11156_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15103__B2 _10601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14997__S _14997_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _19551_/CLK _18997_/D vssd1 vssd1 vccd1 vccd1 _18997_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16778__A _16845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _17948_/A _17954_/C vssd1 vssd1 vccd1 vccd1 _17948_/Y sky130_fd_sc_hd__nor2_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_173_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19659_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_72_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10023__S0 _09782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09964__S0 _09872_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17879_ _17878_/Y _11997_/X _11991_/Y _11998_/Y _12802_/X vssd1 vssd1 vccd1 vccd1
+ _19740_/D sky130_fd_sc_hd__a221oi_1
XFILLER_26_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11715__A _11821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19618_ _19618_/CLK _19618_/D vssd1 vssd1 vccd1 vccd1 _19618_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13417__A1 _19689_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09716__S0 _09793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_188_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19707_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19549_ _19549_/CLK _19549_/D vssd1 vssd1 vccd1 vccd1 _19549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15621__S _15625_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09302_ _14572_/A _18533_/Q _15412_/B _13523_/B _09301_/Y vssd1 vssd1 vccd1 vccd1
+ _09303_/D sky130_fd_sc_hd__o221a_1
XFILLER_80_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09233_ _09854_/A _09233_/B _09233_/C vssd1 vssd1 vccd1 vccd1 _09233_/X sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_111_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19856_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09164_ _18617_/Q _19306_/Q _09190_/A vssd1 vssd1 vccd1 vccd1 _09165_/B sky130_fd_sc_hd__mux2_1
XFILLER_148_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09095_ _18566_/Q vssd1 vssd1 vccd1 vccd1 _11337_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_79_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_126_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _18519_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_163_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17619__A0 _19662_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12156__A1 _14178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13377__A _18376_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09997_ _18839_/Q _19393_/Q _19555_/Q _18807_/Q _09983_/X _09984_/X vssd1 vssd1 vccd1
+ vccd1 _09998_/B sky130_fd_sc_hd__mux4_1
XFILLER_88_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17283__S _17291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15592__A _16992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10014__S0 _09782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10910_ _10910_/A vssd1 vssd1 vccd1 vccd1 _10910_/X sky130_fd_sc_hd__buf_4
XFILLER_45_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12220__S _13529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11890_ _11887_/X _11889_/Y _11801_/A vssd1 vssd1 vccd1 vccd1 _11890_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_71_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10841_ _10837_/Y _10839_/X _10840_/X _10850_/A _10774_/X vssd1 vssd1 vccd1 vccd1
+ _10846_/B sky130_fd_sc_hd__o221a_1
XFILLER_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09627__A3 _09623_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ _13560_/A _13560_/B vssd1 vssd1 vccd1 vccd1 _13561_/A sky130_fd_sc_hd__and2_1
X_10772_ _10772_/A vssd1 vssd1 vccd1 vccd1 _10772_/X sky130_fd_sc_hd__buf_4
XFILLER_44_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12511_ _12511_/A _13711_/A vssd1 vssd1 vccd1 vccd1 _12511_/Y sky130_fd_sc_hd__nor2_4
X_13491_ _18404_/Q _13334_/X _13497_/S vssd1 vssd1 vccd1 vccd1 _13492_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15230_ _18679_/Q _15229_/X _15233_/S vssd1 vssd1 vccd1 vccd1 _15231_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12442_ _12430_/A _12426_/X _12430_/B _12427_/A vssd1 vssd1 vccd1 vccd1 _12450_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_100_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12395__A1 _19756_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15161_ _15161_/A vssd1 vssd1 vccd1 vccd1 _18657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12373_ _12353_/A _14289_/B _12330_/A _14272_/B vssd1 vssd1 vccd1 vccd1 _12373_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_166_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14112_ _14142_/A _14107_/X _14111_/X _13864_/A vssd1 vssd1 vccd1 vccd1 _14112_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09765__A _10011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11324_ _18579_/Q vssd1 vssd1 vccd1 vccd1 _14575_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_126_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15092_ _14559_/A _10834_/X _15092_/S vssd1 vssd1 vccd1 vccd1 _15092_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12147__A1 _19677_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13344__B1 _13338_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18920_ _19442_/CLK _18920_/D vssd1 vssd1 vccd1 vccd1 _18920_/Q sky130_fd_sc_hd__dfxtp_1
X_14043_ _14045_/A _14045_/B vssd1 vssd1 vccd1 vccd1 _14043_/Y sky130_fd_sc_hd__nand2_1
X_11255_ _09756_/B _11224_/Y _11249_/A _11251_/Y _11254_/X vssd1 vssd1 vccd1 vccd1
+ _11255_/X sky130_fd_sc_hd__a221o_1
XFILLER_79_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10206_ _11168_/A _10206_/B vssd1 vssd1 vccd1 vccd1 _10206_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_90_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19861_/CLK sky130_fd_sc_hd__clkbuf_16
X_18851_ _18853_/CLK _18851_/D vssd1 vssd1 vccd1 vccd1 _18851_/Q sky130_fd_sc_hd__dfxtp_1
X_11186_ _18877_/Q _19335_/Q _11186_/S vssd1 vssd1 vccd1 vccd1 _11187_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17802_ _17802_/A vssd1 vssd1 vccd1 vccd1 _19703_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15706__S _15708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10137_ _10140_/A _10134_/X _10136_/X vssd1 vssd1 vccd1 vccd1 _10137_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_39_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13647__A1 _12401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18782_ _19592_/CLK _18782_/D vssd1 vssd1 vccd1 vccd1 _18782_/Q sky130_fd_sc_hd__dfxtp_1
X_15994_ _14879_/X _18996_/Q _15994_/S vssd1 vssd1 vccd1 vccd1 _15995_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17733_ _17737_/A _17737_/C vssd1 vssd1 vccd1 vccd1 _17733_/Y sky130_fd_sc_hd__xnor2_1
X_10068_ _10068_/A _10068_/B vssd1 vssd1 vccd1 vccd1 _10068_/X sky130_fd_sc_hd__or2_1
XFILLER_94_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14945_ _14943_/X _14945_/B _14945_/C vssd1 vssd1 vccd1 vccd1 _14945_/X sky130_fd_sc_hd__and3b_1
XFILLER_48_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17664_ _12713_/X _17662_/Y _17686_/S vssd1 vssd1 vccd1 vccd1 _17664_/X sky130_fd_sc_hd__mux2_1
X_14876_ _14894_/C _14872_/Y _14874_/Y _14875_/X _14842_/X vssd1 vssd1 vccd1 vccd1
+ _14877_/B sky130_fd_sc_hd__o221a_2
XFILLER_165_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19403_ _19597_/CLK _19403_/D vssd1 vssd1 vccd1 vccd1 _19403_/Q sky130_fd_sc_hd__dfxtp_1
X_16615_ _19263_/Q vssd1 vssd1 vccd1 vccd1 _16616_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13827_ _14070_/A vssd1 vssd1 vccd1 vccd1 _13827_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17595_ _19655_/Q _16829_/A _17601_/S vssd1 vssd1 vccd1 vccd1 _17596_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14846__A _16677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10308__S1 _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19334_ _19643_/CLK _19334_/D vssd1 vssd1 vccd1 vccd1 _19334_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12083__A0 _10299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13758_ _13689_/X _13685_/X _13758_/S vssd1 vssd1 vccd1 vccd1 _13758_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16546_ _16546_/A vssd1 vssd1 vccd1 vccd1 _19229_/D sky130_fd_sc_hd__clkbuf_1
X_12709_ _18239_/B _12651_/X _12528_/X _19835_/Q _12708_/X vssd1 vssd1 vccd1 vccd1
+ _12709_/X sky130_fd_sc_hd__a221o_2
X_19265_ _19717_/CLK _19265_/D vssd1 vssd1 vccd1 vccd1 _19265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16477_ _16488_/A vssd1 vssd1 vccd1 vccd1 _16486_/S sky130_fd_sc_hd__buf_4
X_13689_ _14176_/B _14111_/A _13689_/S vssd1 vssd1 vccd1 vccd1 _13689_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18216_ _19859_/Q _18212_/B _18215_/Y vssd1 vssd1 vccd1 vccd1 _19859_/D sky130_fd_sc_hd__o21a_1
X_15428_ _15485_/S vssd1 vssd1 vccd1 vccd1 _15437_/S sky130_fd_sc_hd__buf_2
XFILLER_31_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_19_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19196_ _19614_/CLK _19196_/D vssd1 vssd1 vccd1 vccd1 _19196_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12085__B _13604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17368__S _17374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_43_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19590_/CLK sky130_fd_sc_hd__clkbuf_16
X_18147_ _19835_/Q _18148_/C _19836_/Q vssd1 vssd1 vccd1 vccd1 _18149_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__15677__A _15734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15359_ _15359_/A vssd1 vssd1 vccd1 vccd1 _18728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18053__A _18077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10397__B1 _09315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18078_ _18199_/A vssd1 vssd1 vccd1 vccd1 _18114_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_117_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09920_ _19426_/Q _19202_/Q _19719_/Q _19170_/Q _09914_/A _09770_/X vssd1 vssd1 vccd1
+ vccd1 _09920_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17892__A _17892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17029_ _17029_/A vssd1 vssd1 vccd1 vccd1 _19418_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10149__B1 _09625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10614__A _11028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_58_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19587_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09851_ _18778_/Q _19007_/Q _18938_/Q _19236_/Q _10010_/S _09841_/A vssd1 vssd1 vccd1
+ vccd1 _09852_/B sky130_fd_sc_hd__mux4_1
XFILLER_112_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _09782_/A vssd1 vssd1 vccd1 vccd1 _09782_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_112_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09937__S0 _09803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15351__S _15351_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13271__C1 _13270_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11180__A _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09216_ _10007_/A vssd1 vssd1 vccd1 vccd1 _09217_/A sky130_fd_sc_hd__buf_2
XFILLER_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17278__S _17280_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09147_ _09147_/A vssd1 vssd1 vccd1 vccd1 _09841_/A sky130_fd_sc_hd__buf_2
XFILLER_108_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11040_ _19597_/Q _19435_/Q _18881_/Q _18651_/Q _10959_/X _10969_/A vssd1 vssd1 vccd1
+ vccd1 _11041_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10235__S0 _10224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10243__B _10243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10786__S1 _10785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16211__A _18207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14826__B1 _14824_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _12991_/A vssd1 vssd1 vccd1 vccd1 _13034_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14730_ _14729_/X _18587_/Q _14762_/S vssd1 vssd1 vccd1 vccd1 _14731_/A sky130_fd_sc_hd__mux2_1
X_11942_ _11511_/A _11470_/A _12024_/A vssd1 vssd1 vccd1 vccd1 _11942_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10459__A1_N _18438_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _14677_/A _17781_/B vssd1 vssd1 vccd1 vccd1 _14662_/A sky130_fd_sc_hd__and2_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _11746_/A _11746_/B _11747_/A _11787_/A _11846_/A vssd1 vssd1 vccd1 vccd1
+ _11873_/X sky130_fd_sc_hd__o2111a_1
XANTENNA__14666__A _14677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ _13769_/S vssd1 vssd1 vccd1 vccd1 _13759_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13570__A _13570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16400_ _19165_/Q _15548_/X _16402_/S vssd1 vssd1 vccd1 vccd1 _16401_/A sky130_fd_sc_hd__mux2_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ _19505_/Q _19119_/Q _19569_/Q _18725_/Q _11027_/S _10813_/A vssd1 vssd1 vccd1
+ vccd1 _10825_/B sky130_fd_sc_hd__mux4_1
XFILLER_60_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17380_ _17380_/A vssd1 vssd1 vccd1 vccd1 _19559_/D sky130_fd_sc_hd__clkbuf_1
X_14592_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14640_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16331_ _16342_/A vssd1 vssd1 vccd1 vccd1 _16340_/S sky130_fd_sc_hd__buf_4
X_13543_ _13543_/A vssd1 vssd1 vccd1 vccd1 _18419_/D sky130_fd_sc_hd__clkbuf_1
X_10755_ _10866_/A _10755_/B vssd1 vssd1 vccd1 vccd1 _10755_/X sky130_fd_sc_hd__or2_1
XFILLER_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16262_ _16103_/X _19104_/Q _16268_/S vssd1 vssd1 vccd1 vccd1 _16263_/A sky130_fd_sc_hd__mux2_1
X_19050_ _19633_/CLK _19050_/D vssd1 vssd1 vccd1 vccd1 _19050_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_20_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13474_ _13474_/A vssd1 vssd1 vccd1 vccd1 _18396_/D sky130_fd_sc_hd__clkbuf_1
X_10686_ _19604_/Q _19442_/Q _18888_/Q _18658_/Q _10860_/S _09139_/A vssd1 vssd1 vccd1
+ vccd1 _10687_/B sky130_fd_sc_hd__mux4_1
XFILLER_173_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15213_ _16715_/A vssd1 vssd1 vccd1 vccd1 _15213_/X sky130_fd_sc_hd__clkbuf_2
X_18001_ _18027_/A _18006_/C vssd1 vssd1 vccd1 vccd1 _18001_/Y sky130_fd_sc_hd__nor2_1
X_12425_ _12426_/A _14324_/B vssd1 vssd1 vccd1 vccd1 _12427_/A sky130_fd_sc_hd__and2_1
X_16193_ _16193_/A vssd1 vssd1 vccd1 vccd1 _19069_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15144_ _18652_/Q _15143_/X _15153_/S vssd1 vssd1 vccd1 vccd1 _15145_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10474__S0 _09631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ _12330_/A _14272_/B _12371_/B _12333_/B vssd1 vssd1 vccd1 vccd1 _12357_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14431__D_N _13529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ _11381_/C _11306_/X input33/X vssd1 vssd1 vccd1 vccd1 _11462_/A sky130_fd_sc_hd__o21ba_2
X_15075_ _16740_/A vssd1 vssd1 vccd1 vccd1 _16844_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16820__S _16823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12287_ _12233_/A _14227_/B _12262_/A _14241_/B vssd1 vssd1 vccd1 vccd1 _12287_/X
+ sky130_fd_sc_hd__o22a_1
X_18903_ _19587_/CLK _18903_/D vssd1 vssd1 vccd1 vccd1 _18903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output74_A _11926_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14026_ _14026_/A _14026_/B vssd1 vssd1 vccd1 vccd1 _14026_/Y sky130_fd_sc_hd__nor2_1
X_11238_ _11238_/A _11238_/B vssd1 vssd1 vccd1 vccd1 _11266_/B sky130_fd_sc_hd__nor2_1
XFILLER_45_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10777__S1 _10713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18834_ _19713_/CLK _18834_/D vssd1 vssd1 vccd1 vccd1 _18834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11169_ _18845_/Q _19399_/Q _19561_/Q _18813_/Q _11153_/X _09542_/A vssd1 vssd1 vccd1
+ vccd1 _11169_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18765_ _19513_/CLK _18765_/D vssd1 vssd1 vccd1 vccd1 _18765_/Q sky130_fd_sc_hd__dfxtp_1
X_15977_ _14782_/X _18988_/Q _15983_/S vssd1 vssd1 vccd1 vccd1 _15978_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09839__A3 _09837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17716_ _17716_/A _17720_/C vssd1 vssd1 vccd1 vccd1 _17716_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_36_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14928_ _16699_/A vssd1 vssd1 vccd1 vccd1 _16803_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18696_ _19636_/CLK _18696_/D vssd1 vssd1 vccd1 vccd1 _18696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17647_ _19667_/Q _17646_/X _17653_/S vssd1 vssd1 vccd1 vccd1 _17648_/A sky130_fd_sc_hd__mux2_1
X_14859_ _14873_/A _14859_/B _14859_/C _14859_/D vssd1 vssd1 vccd1 vccd1 _14859_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17578_ _17578_/A vssd1 vssd1 vccd1 vccd1 _19647_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19317_ _19543_/CLK _19317_/D vssd1 vssd1 vccd1 vccd1 _19317_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10606__A1 _09169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16529_ _16529_/A vssd1 vssd1 vccd1 vccd1 _19221_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10609__A _10956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19248_ _19634_/CLK _19248_/D vssd1 vssd1 vccd1 vccd1 _19248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19179_ _19630_/CLK _19179_/D vssd1 vssd1 vccd1 vccd1 _19179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15200__A _16702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09903_ _09919_/A _09903_/B vssd1 vssd1 vccd1 vccd1 _09903_/X sky130_fd_sc_hd__or2_1
XANTENNA__14520__A2 _12692_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09834_ _19427_/Q _19203_/Q _19720_/Q _19171_/Q _09874_/S _09810_/A vssd1 vssd1 vccd1
+ vccd1 _09834_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _10011_/S vssd1 vssd1 vccd1 vccd1 _10010_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_101_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16966__A _16977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09386__S1 _09364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09696_ _09704_/A vssd1 vssd1 vccd1 vccd1 _09697_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17222__A1 _12779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16177__S _16183_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12718__B _18631_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16905__S _16913_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ _18596_/Q _19285_/Q _10540_/S vssd1 vssd1 vccd1 vccd1 _10540_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10471_ _11102_/A _10471_/B vssd1 vssd1 vccd1 vccd1 _10471_/X sky130_fd_sc_hd__or2_1
XFILLER_41_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12210_ _12210_/A _12237_/A vssd1 vssd1 vccd1 vccd1 _12235_/A sky130_fd_sc_hd__or2_2
X_13190_ _19664_/Q _12737_/A _13205_/A _18388_/Q vssd1 vssd1 vccd1 vccd1 _13190_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12453__B _13529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12141_ _12141_/A _12141_/B vssd1 vssd1 vccd1 vccd1 _12142_/A sky130_fd_sc_hd__xnor2_4
XFILLER_68_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12072_ _12072_/A vssd1 vssd1 vccd1 vccd1 _12072_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10759__S1 _09353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ _09925_/A _11012_/X _11021_/X _09305_/A _11022_/X vssd1 vssd1 vccd1 vccd1
+ _12460_/A sky130_fd_sc_hd__a32o_4
X_15900_ _14808_/X _18953_/Q _15902_/S vssd1 vssd1 vccd1 vccd1 _15901_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13565__A _15095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16880_ _19353_/Q _16686_/X _16880_/S vssd1 vssd1 vccd1 vccd1 _16881_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13284__B _18633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15831_ _15831_/A vssd1 vssd1 vccd1 vccd1 _18922_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18550_ _19481_/CLK _18550_/D vssd1 vssd1 vccd1 vccd1 _18550_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ _18303_/Q _18304_/Q _18306_/Q _18305_/Q vssd1 vssd1 vccd1 vccd1 _12984_/D
+ sky130_fd_sc_hd__and4_1
X_15762_ _15762_/A vssd1 vssd1 vccd1 vccd1 _18891_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17501_ _19613_/Q _16693_/X _17507_/S vssd1 vssd1 vccd1 vccd1 _17502_/A sky130_fd_sc_hd__mux2_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ _16639_/A vssd1 vssd1 vccd1 vccd1 _16743_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ _11925_/A _11925_/B vssd1 vssd1 vccd1 vccd1 _11930_/B sky130_fd_sc_hd__xnor2_4
XFILLER_61_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18481_ _18482_/CLK _18481_/D vssd1 vssd1 vccd1 vccd1 _18481_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _18861_/Q _15529_/X _15697_/S vssd1 vssd1 vccd1 vccd1 _15694_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _17432_/A vssd1 vssd1 vccd1 vccd1 _19582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11856_ _18357_/Q vssd1 vssd1 vccd1 vccd1 _13215_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14644_ input39/X _14640_/X _14643_/X _14547_/A vssd1 vssd1 vccd1 vccd1 _14645_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10049__C1 _09395_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ _10807_/A _10807_/B vssd1 vssd1 vccd1 vccd1 _10807_/X sky130_fd_sc_hd__or2_1
X_17363_ _16806_/X _19552_/Q _17363_/S vssd1 vssd1 vccd1 vccd1 _17364_/A sky130_fd_sc_hd__mux2_1
X_14575_ _14575_/A _14580_/B vssd1 vssd1 vccd1 vccd1 _14575_/X sky130_fd_sc_hd__or2_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11787_ _11787_/A _11787_/B vssd1 vssd1 vccd1 vccd1 _11787_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19102_ _19616_/CLK _19102_/D vssd1 vssd1 vccd1 vccd1 _19102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16314_ _16074_/X _19127_/Q _16318_/S vssd1 vssd1 vccd1 vccd1 _16315_/A sky130_fd_sc_hd__mux2_1
X_10738_ _10858_/A _18855_/Q vssd1 vssd1 vccd1 vccd1 _10738_/Y sky130_fd_sc_hd__nor2_1
X_13526_ _13526_/A _13526_/B _13526_/C vssd1 vssd1 vccd1 vccd1 _13545_/B sky130_fd_sc_hd__or3_2
X_17294_ _19521_/Q _16705_/X _17302_/S vssd1 vssd1 vccd1 vccd1 _17295_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19033_ _19648_/CLK _19033_/D vssd1 vssd1 vccd1 vccd1 _19033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13457_ _13457_/A vssd1 vssd1 vccd1 vccd1 _18388_/D sky130_fd_sc_hd__clkbuf_1
X_16245_ _16245_/A vssd1 vssd1 vccd1 vccd1 _19096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10669_ _10669_/A _18856_/Q vssd1 vssd1 vccd1 vccd1 _10669_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14637__A1_N input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12408_ _12408_/A _12408_/B vssd1 vssd1 vccd1 vccd1 _12408_/Y sky130_fd_sc_hd__nor2_1
X_13388_ _13388_/A _13413_/B vssd1 vssd1 vccd1 vccd1 _13388_/X sky130_fd_sc_hd__or2_1
X_16176_ _16176_/A vssd1 vssd1 vccd1 vccd1 _19061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12363__B _14284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput106 _09109_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_ld_type[1] sky130_fd_sc_hd__buf_2
XFILLER_99_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput117 _12483_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[15] sky130_fd_sc_hd__buf_2
X_12339_ _11980_/X _12337_/X _12338_/X _12193_/X vssd1 vssd1 vccd1 vccd1 _12339_/X
+ sky130_fd_sc_hd__o211a_1
X_15127_ _18645_/Q _15123_/X _15125_/X _11222_/A vssd1 vssd1 vccd1 vccd1 _18645_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15955__A _15955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput128 _12499_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[25] sky130_fd_sc_hd__buf_2
XANTENNA__16550__S _16558_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput139 _12468_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[6] sky130_fd_sc_hd__buf_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18229__B1 _12948_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15058_ _18488_/Q _15059_/B vssd1 vssd1 vccd1 vccd1 _15069_/B sky130_fd_sc_hd__nand2_1
XFILLER_141_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14009_ _14005_/B _13658_/X _13863_/A _14008_/X vssd1 vssd1 vccd1 vccd1 _14009_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19866_ _19866_/CLK _19866_/D vssd1 vssd1 vccd1 vccd1 _19866_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09164__S _09190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18817_ _18982_/CLK _18817_/D vssd1 vssd1 vccd1 vccd1 _18817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19797_ _19798_/CLK _19797_/D vssd1 vssd1 vccd1 vccd1 _19797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17381__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09550_ _10475_/A vssd1 vssd1 vccd1 vccd1 _10432_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18748_ _19592_/CLK _18748_/D vssd1 vssd1 vccd1 vccd1 _18748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09481_ _09481_/A vssd1 vssd1 vccd1 vccd1 _09482_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18679_ _19625_/CLK _18679_/D vssd1 vssd1 vccd1 vccd1 _18679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11723__A _11723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16460__S _16464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09817_ _09806_/Y _09812_/Y _09814_/Y _09816_/Y _09940_/A vssd1 vssd1 vccd1 vccd1
+ _09817_/X sky130_fd_sc_hd__o221a_2
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16696__A _16696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17291__S _17291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15804__S _15806_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ _19623_/Q _19461_/Q _18907_/Q _18677_/Q _09734_/X _10186_/A vssd1 vssd1 vccd1
+ vccd1 _09748_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _09679_/A vssd1 vssd1 vccd1 vccd1 _11123_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09684__A1 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11710_ _12017_/B vssd1 vssd1 vccd1 vccd1 _12390_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__10913__S1 _10910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _13442_/C vssd1 vssd1 vccd1 vccd1 _13536_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11641_ _11343_/X _11640_/Y _11584_/A _11357_/Y vssd1 vssd1 vccd1 vccd1 _11643_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17320__A _17376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14360_ _14360_/A vssd1 vssd1 vccd1 vccd1 _18464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11572_ _11572_/A vssd1 vssd1 vccd1 vccd1 _11572_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17903__C1 _12802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13311_ _13311_/A vssd1 vssd1 vccd1 vccd1 _13311_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10523_ _19607_/Q _19445_/Q _18891_/Q _18661_/Q _10500_/X _10238_/A vssd1 vssd1 vccd1
+ vccd1 _10524_/B sky130_fd_sc_hd__mux4_2
Xinput19 io_dbus_rdata[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_2
XFILLER_167_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14291_ _13795_/X _14286_/X _14288_/Y _14290_/X vssd1 vssd1 vccd1 vccd1 _14291_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__12464__A _12464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13242_ _18312_/Q _13130_/X _12749_/X _19801_/Q vssd1 vssd1 vccd1 vccd1 _13242_/X
+ sky130_fd_sc_hd__a22o_1
X_16030_ _16030_/A vssd1 vssd1 vccd1 vccd1 _19012_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10429__S0 _09632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10454_ _19415_/Q _19191_/Q _19708_/Q _19159_/Q _10401_/A _10245_/A vssd1 vssd1 vccd1
+ vccd1 _10454_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17466__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ _18354_/Q _13115_/A _12671_/A _18683_/Q _13172_/X vssd1 vssd1 vccd1 vccd1
+ _13173_/X sky130_fd_sc_hd__a221o_1
X_10385_ _19257_/Q _19028_/Q _18959_/Q _19353_/Q _10277_/S _10384_/X vssd1 vssd1 vccd1
+ vccd1 _10386_/B sky130_fd_sc_hd__mux4_1
XFILLER_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12124_ _12091_/A _12122_/Y _12169_/C _11859_/X vssd1 vssd1 vccd1 vccd1 _12124_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_124_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17981_ _19779_/Q _17981_/B vssd1 vssd1 vccd1 vccd1 _17988_/C sky130_fd_sc_hd__and2_2
XFILLER_124_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13299__A2 _12603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14496__A1 _19756_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19720_ _19720_/CLK _19720_/D vssd1 vssd1 vccd1 vccd1 _19720_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13295__A _13295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11808__A _13984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16932_ _16932_/A vssd1 vssd1 vccd1 vccd1 _19375_/D sky130_fd_sc_hd__clkbuf_1
X_12055_ _12155_/A _12055_/B vssd1 vssd1 vccd1 vccd1 _12131_/C sky130_fd_sc_hd__nand2_1
XANTENNA__10712__A _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11006_ _19244_/Q _19015_/Q _18946_/Q _19340_/Q _10724_/A _10712_/A vssd1 vssd1 vccd1
+ vccd1 _11006_/X sky130_fd_sc_hd__mux4_2
X_19651_ _19838_/CLK _19651_/D vssd1 vssd1 vccd1 vccd1 _19651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16863_ _19345_/Q _16661_/X _16869_/S vssd1 vssd1 vccd1 vccd1 _16864_/A sky130_fd_sc_hd__mux2_1
X_18602_ _19581_/CLK _18602_/D vssd1 vssd1 vccd1 vccd1 _18602_/Q sky130_fd_sc_hd__dfxtp_1
X_15814_ _15814_/A vssd1 vssd1 vccd1 vccd1 _18914_/D sky130_fd_sc_hd__clkbuf_1
X_19582_ _19712_/CLK _19582_/D vssd1 vssd1 vccd1 vccd1 _19582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16794_ _16826_/A vssd1 vssd1 vccd1 vccd1 _16807_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18533_ _18548_/CLK _18533_/D vssd1 vssd1 vccd1 vccd1 _18533_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17198__A0 _18443_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15745_ _14753_/X _18884_/Q _15747_/S vssd1 vssd1 vccd1 vccd1 _15746_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12957_ _18296_/Q _18295_/Q _12957_/C vssd1 vssd1 vccd1 vccd1 _12959_/B sky130_fd_sc_hd__and3_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11908_ _13246_/A _11962_/D vssd1 vssd1 vccd1 vccd1 _11936_/B sky130_fd_sc_hd__nand2_1
X_18464_ _18471_/CLK _18464_/D vssd1 vssd1 vccd1 vccd1 _18464_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15676_ _15676_/A vssd1 vssd1 vccd1 vccd1 _18853_/D sky130_fd_sc_hd__clkbuf_1
X_12888_ _18275_/Q _12884_/C _12887_/Y vssd1 vssd1 vccd1 vccd1 _18275_/D sky130_fd_sc_hd__o21a_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _17461_/S vssd1 vssd1 vccd1 vccd1 _17424_/S sky130_fd_sc_hd__buf_6
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14627_ _18563_/Q _14613_/X _14622_/X input65/X vssd1 vssd1 vccd1 vccd1 _14628_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10690__C1 _09244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18395_ _18395_/CLK _18395_/D vssd1 vssd1 vccd1 vccd1 _18395_/Q sky130_fd_sc_hd__dfxtp_1
X_11839_ _11939_/A _11839_/B vssd1 vssd1 vccd1 vccd1 _11842_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__16545__S _16547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10159__A _10212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17346_ _16781_/X _19544_/Q _17352_/S vssd1 vssd1 vccd1 vccd1 _17347_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14558_ _18540_/Q _14550_/X _14557_/X _14548_/X vssd1 vssd1 vccd1 vccd1 _18540_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13509_ _13509_/A vssd1 vssd1 vccd1 vccd1 _18412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17277_ _17277_/A vssd1 vssd1 vccd1 vccd1 _19513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14489_ _14591_/B vssd1 vssd1 vccd1 vccd1 _14498_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_9_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19016_ _19633_/CLK _19016_/D vssd1 vssd1 vccd1 vccd1 _19016_/Q sky130_fd_sc_hd__dfxtp_1
X_16228_ _16228_/A vssd1 vssd1 vccd1 vccd1 _19088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16159_ _16061_/X _19054_/Q _16161_/S vssd1 vssd1 vccd1 vccd1 _16160_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18061__A _18077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10840__S0 _10711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14487__A1 _19752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10622__A _10622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_142_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19849_ _19851_/CLK _19849_/D vssd1 vssd1 vccd1 vccd1 _19849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09602_ _09602_/A vssd1 vssd1 vccd1 vccd1 _09603_/A sky130_fd_sc_hd__buf_2
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09533_ _18456_/Q _09308_/A _09428_/A _09532_/X vssd1 vssd1 vccd1 vccd1 _12504_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_58_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11453__A input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16936__A0 _16765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ _19531_/Q _19145_/Q _19595_/Q _18751_/Q _10350_/S _09442_/X vssd1 vssd1 vccd1
+ vccd1 _09465_/B sky130_fd_sc_hd__mux4_1
XFILLER_58_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10681__C1 _10823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09395_ _09395_/A vssd1 vssd1 vccd1 vccd1 _09395_/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__13214__A2 _13212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17140__A _17245_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_67_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10984__B1 _09177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13099__B _13104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16190__S _16194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10831__S0 _09152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10170_ _10163_/X _10165_/X _10167_/X _10169_/X _09249_/A vssd1 vssd1 vccd1 vccd1
+ _10170_/X sky130_fd_sc_hd__a221o_1
XFILLER_161_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11433__A2_N _18417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14939__A _16702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13860_ _14092_/A vssd1 vssd1 vccd1 vccd1 _14323_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09532__S _10494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12811_ _18034_/A vssd1 vssd1 vccd1 vccd1 _18225_/A sky130_fd_sc_hd__buf_4
XANTENNA__12459__A _12459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13791_ _13880_/S vssd1 vssd1 vccd1 vccd1 _13888_/S sky130_fd_sc_hd__buf_2
XANTENNA__14650__A1 _14553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09657__B2 _18453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14650__B2 input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15530_ _18797_/Q _15529_/X _15536_/S vssd1 vssd1 vccd1 vccd1 _15531_/A sky130_fd_sc_hd__mux2_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12742_ _12742_/A vssd1 vssd1 vccd1 vccd1 _13154_/B sky130_fd_sc_hd__buf_2
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10898__S0 _10648_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16927__A0 _16752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11082__B _11082_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12673_ _18382_/Q _12568_/X _12642_/A _18353_/Q vssd1 vssd1 vccd1 vccd1 _12673_/X
+ sky130_fd_sc_hd__a22o_1
X_15461_ _15472_/A vssd1 vssd1 vccd1 vccd1 _15470_/S sky130_fd_sc_hd__buf_4
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16365__S _16369_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _17200_/A vssd1 vssd1 vccd1 vccd1 _19486_/D sky130_fd_sc_hd__clkbuf_1
X_14412_ _14426_/A vssd1 vssd1 vccd1 vccd1 _14424_/S sky130_fd_sc_hd__clkbuf_2
X_11624_ _11624_/A _11624_/B vssd1 vssd1 vccd1 vccd1 _11624_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18180_ _19847_/Q _18183_/C _18170_/X vssd1 vssd1 vccd1 vccd1 _18180_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09768__A _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15392_ _15392_/A vssd1 vssd1 vccd1 vccd1 _18743_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15489__B _15592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17131_ _17131_/A vssd1 vssd1 vccd1 vccd1 _19464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11810__B _11843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17352__A0 _16790_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14343_ _18459_/Q _18491_/Q _14352_/S vssd1 vssd1 vccd1 vccd1 _14344_/A sky130_fd_sc_hd__mux2_1
X_11555_ _11314_/A _11599_/A vssd1 vssd1 vccd1 vccd1 _11556_/A sky130_fd_sc_hd__and2b_1
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10506_ _09927_/X _10494_/X _10505_/X _09307_/A _18437_/Q vssd1 vssd1 vccd1 vccd1
+ _12478_/B sky130_fd_sc_hd__a32o_4
X_14274_ _14274_/A _14274_/B vssd1 vssd1 vccd1 vccd1 _14274_/X sky130_fd_sc_hd__or2_1
X_17062_ _19434_/Q _16740_/X _17062_/S vssd1 vssd1 vccd1 vccd1 _17063_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12302__A1_N _14575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11486_ _11282_/A _14543_/A _11550_/B _11474_/A vssd1 vssd1 vccd1 vccd1 _13977_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12716__A1 _13106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16013_ _16013_/A vssd1 vssd1 vccd1 vccd1 _19004_/D sky130_fd_sc_hd__clkbuf_1
X_13225_ _17954_/B _12629_/S _13224_/X vssd1 vssd1 vccd1 vccd1 _13225_/X sky130_fd_sc_hd__o21a_1
X_10437_ _18829_/Q _19383_/Q _19545_/Q _18797_/Q _11112_/S _10384_/X vssd1 vssd1 vccd1
+ vccd1 _10438_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13156_ _13156_/A vssd1 vssd1 vccd1 vccd1 _13326_/B sky130_fd_sc_hd__clkbuf_2
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _10368_/A vssd1 vssd1 vccd1 vccd1 _10368_/X sky130_fd_sc_hd__buf_2
XFILLER_152_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _12155_/A _12079_/B _12081_/B _13567_/A vssd1 vssd1 vccd1 vccd1 _12108_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_3_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17964_ _17980_/A _17964_/B _17965_/B vssd1 vssd1 vccd1 vccd1 _19772_/D sky130_fd_sc_hd__nor3_1
X_13087_ _13297_/A _13076_/Y _13086_/X _13306_/A _18626_/Q vssd1 vssd1 vccd1 vccd1
+ _13088_/A sky130_fd_sc_hd__a32o_2
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15130__A2 _13873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10299_ _10299_/A _12485_/A vssd1 vssd1 vccd1 vccd1 _10300_/B sky130_fd_sc_hd__nor2_1
X_19703_ _19703_/CLK _19703_/D vssd1 vssd1 vccd1 vccd1 _19703_/Q sky130_fd_sc_hd__dfxtp_1
X_12038_ _12010_/A _13595_/A _12037_/X vssd1 vssd1 vccd1 vccd1 _12038_/X sky130_fd_sc_hd__o21a_1
X_16915_ _19369_/Q _16737_/X _16917_/S vssd1 vssd1 vccd1 vccd1 _16916_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17895_ _17895_/A vssd1 vssd1 vccd1 vccd1 _17895_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09896__B2 _09895_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15444__S _15448_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19634_ _19634_/CLK _19634_/D vssd1 vssd1 vccd1 vccd1 _19634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16846_ _16846_/A vssd1 vssd1 vccd1 vccd1 _19338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09991__S1 _09984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19565_ _19598_/CLK _19565_/D vssd1 vssd1 vccd1 vccd1 _19565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16777_ _16777_/A vssd1 vssd1 vccd1 vccd1 _16777_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13989_ _11813_/Y _13827_/X _13988_/X _13828_/X vssd1 vssd1 vccd1 vccd1 _13989_/X
+ sky130_fd_sc_hd__a211o_1
X_18516_ _18519_/CLK _18516_/D vssd1 vssd1 vccd1 vccd1 _18516_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15728_ _18877_/Q _15580_/X _15730_/S vssd1 vssd1 vccd1 vccd1 _15729_/A sky130_fd_sc_hd__mux2_1
X_19496_ _19496_/CLK _19496_/D vssd1 vssd1 vccd1 vccd1 _19496_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10889__S0 _10711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18447_ _19468_/CLK _18447_/D vssd1 vssd1 vccd1 vccd1 _18447_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16275__S _16279_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15659_ _15659_/A vssd1 vssd1 vccd1 vccd1 _18846_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14584__A _14584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09180_ _09451_/A vssd1 vssd1 vccd1 vccd1 _09549_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18378_ _19690_/CLK _18378_/D vssd1 vssd1 vccd1 vccd1 _18378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12955__A1 _18295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11720__B _11720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17895__A _17895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17329_ _17329_/A vssd1 vssd1 vccd1 vccd1 _19536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12707__A1 _19670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15619__S _15625_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13380__A1 _18294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17646__A1 _17645_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17834__S _17838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15121__A2 _15116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10782__A1_N _18432_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15354__S _15362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09516_ _19433_/Q _19209_/Q _19726_/Q _19177_/Q _10450_/S _09587_/A vssd1 vssd1 vccd1
+ vccd1 _09516_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09447_ _09447_/A vssd1 vssd1 vccd1 vccd1 _09448_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11911__A _14587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09588__A _10451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09378_ _10593_/A vssd1 vssd1 vccd1 vccd1 _10395_/A sky130_fd_sc_hd__buf_2
XFILLER_71_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12726__B _12726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16913__S _16913_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11340_ _11285_/A _11528_/B _11339_/X vssd1 vssd1 vccd1 vccd1 _11477_/A sky130_fd_sc_hd__o21ai_1
XFILLER_153_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11271_ _11271_/A _11271_/B vssd1 vssd1 vccd1 vccd1 _11274_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12742__A _12742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ _18316_/Q vssd1 vssd1 vccd1 vccd1 _13015_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13371__A1 _12840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10222_ _10447_/A _10222_/B vssd1 vssd1 vccd1 vccd1 _10222_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10804__S0 _10724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ _18604_/Q _19293_/Q _10153_/S vssd1 vssd1 vccd1 vccd1 _10153_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10262__A _10262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11077__B _12473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input36_A io_ibus_inst[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ _10007_/X _10074_/X _10078_/X _10083_/X _09135_/A vssd1 vssd1 vccd1 vccd1
+ _10084_/X sky130_fd_sc_hd__a311o_1
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14961_ input14/X _14960_/X _14925_/X vssd1 vssd1 vccd1 vccd1 _14961_/X sky130_fd_sc_hd__a21o_1
XFILLER_48_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14669__A _14677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16700_ _19293_/Q _16699_/X _16703_/S vssd1 vssd1 vccd1 vccd1 _16701_/A sky130_fd_sc_hd__mux2_1
X_13912_ _18429_/Q _13736_/X _13910_/X _13911_/X vssd1 vssd1 vccd1 vccd1 _18429_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_87_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17680_ _13294_/X _17679_/Y _17686_/S vssd1 vssd1 vccd1 vccd1 _17680_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14892_ _14892_/A vssd1 vssd1 vccd1 vccd1 _18601_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16631_ _19271_/Q vssd1 vssd1 vccd1 vccd1 _16632_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13843_ _13619_/X _13638_/X _13880_/S vssd1 vssd1 vccd1 vccd1 _13843_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10893__C1 _09391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14623__A1 _18562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19350_ _19610_/CLK _19350_/D vssd1 vssd1 vccd1 vccd1 _19350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16562_ _16562_/A vssd1 vssd1 vccd1 vccd1 _19236_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10201__S _10256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13774_ _13742_/S _13720_/A _13996_/B vssd1 vssd1 vccd1 vccd1 _13774_/Y sky130_fd_sc_hd__a21boi_1
X_10986_ _18754_/Q _18983_/Q _18914_/Q _19212_/Q _10668_/A _10906_/A vssd1 vssd1 vccd1
+ vccd1 _10986_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18301_ _19856_/CLK _18301_/D vssd1 vssd1 vccd1 vccd1 _18301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15513_ _16768_/A vssd1 vssd1 vccd1 vccd1 _15513_/X sky130_fd_sc_hd__buf_2
X_12725_ _19804_/Q _12665_/X _12602_/X _18315_/Q _12724_/X vssd1 vssd1 vccd1 vccd1
+ _12726_/B sky130_fd_sc_hd__a221o_2
X_19281_ _19571_/CLK _19281_/D vssd1 vssd1 vccd1 vccd1 _19281_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16376__A1 _15513_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16493_ _16122_/X _19206_/Q _16497_/S vssd1 vssd1 vccd1 vccd1 _16494_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12917__A _12991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18232_ _18250_/A _18232_/B vssd1 vssd1 vccd1 vccd1 _18232_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11821__A _11821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09498__A _10650_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15444_ _18765_/Q _15178_/X _15448_/S vssd1 vssd1 vccd1 vccd1 _15445_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12656_ _13092_/S _12656_/B vssd1 vssd1 vccd1 vccd1 _12656_/X sky130_fd_sc_hd__and2b_1
XFILLER_129_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12937__A1 _18289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18163_ _19841_/Q _18164_/C _19842_/Q vssd1 vssd1 vccd1 vccd1 _18165_/B sky130_fd_sc_hd__a21oi_1
XFILLER_157_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11607_ _11372_/A _11347_/Y _11602_/Y _11604_/X _11606_/X vssd1 vssd1 vccd1 vccd1
+ _11686_/D sky130_fd_sc_hd__a2111oi_4
X_12587_ _12587_/A vssd1 vssd1 vccd1 vccd1 _12674_/A sky130_fd_sc_hd__buf_2
XFILLER_129_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15375_ _15397_/A vssd1 vssd1 vccd1 vccd1 _15384_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16823__S _16823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10948__B1 _10774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17114_ _17114_/A vssd1 vssd1 vccd1 vccd1 _19456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14326_ _13795_/X _14321_/X _14323_/Y _14325_/X vssd1 vssd1 vccd1 vccd1 _14326_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_157_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18094_ _18094_/A _19818_/Q _18094_/C vssd1 vssd1 vccd1 vccd1 _18096_/B sky130_fd_sc_hd__and3_1
XFILLER_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11538_ _11538_/A _11538_/B _11538_/C _11538_/D vssd1 vssd1 vccd1 vccd1 _11538_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_144_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17045_ _19426_/Q _16715_/X _17047_/S vssd1 vssd1 vccd1 vccd1 _17046_/A sky130_fd_sc_hd__mux2_1
X_14257_ _13823_/A _14002_/X _14256_/X _14115_/X vssd1 vssd1 vccd1 vccd1 _14257_/X
+ sky130_fd_sc_hd__a211o_1
X_11469_ _11966_/B vssd1 vssd1 vccd1 vccd1 _12344_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_171_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17628__A1 _17627_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13208_ _18309_/Q _13130_/A _12582_/A _19862_/Q vssd1 vssd1 vccd1 vccd1 _13208_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14188_ _14192_/A _14192_/B vssd1 vssd1 vccd1 vccd1 _14188_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15963__A _16031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13139_ _13311_/A vssd1 vssd1 vccd1 vccd1 _13139_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18996_ _19223_/CLK _18996_/D vssd1 vssd1 vccd1 vccd1 _18996_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10271__S1 _09145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17947_ _17957_/D vssd1 vssd1 vccd1 vccd1 _17954_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11125__B1 _09681_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_15_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10023__S1 _09979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__S1 _09869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17878_ _17878_/A vssd1 vssd1 vccd1 vccd1 _17878_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19617_ _19716_/CLK _19617_/D vssd1 vssd1 vccd1 vccd1 _19617_/Q sky130_fd_sc_hd__dfxtp_1
X_16829_ _16829_/A vssd1 vssd1 vccd1 vccd1 _16829_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13417__A2 _12703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15811__A0 _14714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15902__S _15902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19548_ _19624_/CLK _19548_/D vssd1 vssd1 vccd1 vccd1 _19548_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09716__S1 _09704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14090__A2 _14093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09301_ _18575_/Q _16212_/A vssd1 vssd1 vccd1 vccd1 _09301_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_55_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19479_ _19488_/CLK _19479_/D vssd1 vssd1 vccd1 vccd1 _19479_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16367__A1 _15500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09232_ _09237_/A _09219_/X _09221_/X _09231_/X vssd1 vssd1 vccd1 vccd1 _09233_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15203__A _16705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09201__A _10313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09163_ _09163_/A vssd1 vssd1 vccd1 vccd1 _09190_/A sky130_fd_sc_hd__buf_2
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10347__A _11135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09094_ _09094_/A vssd1 vssd1 vccd1 vccd1 _12495_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_162_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13658__A _13658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15349__S _15351_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16034__A _16847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13353__A1 _12779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11178__A _11178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17564__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10082__A _10212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09996_ _09996_/A vssd1 vssd1 vccd1 vccd1 _10020_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15592__B _15592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14489__A _14591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14853__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10014__S1 _09979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10840_ _19248_/Q _19019_/Q _18950_/Q _19344_/Q _10711_/A _10713_/X vssd1 vssd1 vccd1
+ vccd1 _10840_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10771_ _10634_/A _10770_/X _10797_/A vssd1 vssd1 vccd1 vccd1 _10771_/X sky130_fd_sc_hd__a21o_1
XFILLER_71_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12510_ _13747_/S _12510_/B vssd1 vssd1 vccd1 vccd1 _13711_/A sky130_fd_sc_hd__nor2_1
X_13490_ _13490_/A vssd1 vssd1 vccd1 vccd1 _18403_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15030__A1 _14744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12441_ _19758_/Q _12186_/X _12437_/X _12440_/X vssd1 vssd1 vccd1 vccd1 _12441_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_139_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12372_ _12372_/A vssd1 vssd1 vccd1 vccd1 _14289_/B sky130_fd_sc_hd__buf_2
X_15160_ _18657_/Q _15159_/X _15169_/S vssd1 vssd1 vccd1 vccd1 _15161_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09891__S0 _09809_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14111_ _14111_/A _12008_/A vssd1 vssd1 vccd1 vccd1 _14111_/X sky130_fd_sc_hd__or2b_1
X_11323_ _18580_/Q vssd1 vssd1 vccd1 vccd1 _14578_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15091_ _15091_/A vssd1 vssd1 vccd1 vccd1 _18622_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12472__A _12472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14042_ _14126_/A _14045_/B _14041_/X vssd1 vssd1 vccd1 vccd1 _14042_/Y sky130_fd_sc_hd__o21ai_1
X_11254_ _11254_/A _11254_/B _11254_/C _11253_/X vssd1 vssd1 vccd1 vccd1 _11254_/X
+ sky130_fd_sc_hd__or4b_2
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17474__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ _18770_/Q _18999_/Q _18930_/Q _19228_/Q _09545_/S _10080_/A vssd1 vssd1 vccd1
+ vccd1 _10206_/B sky130_fd_sc_hd__mux4_1
XFILLER_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18850_ _19534_/CLK _18850_/D vssd1 vssd1 vccd1 vccd1 _18850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11185_ _11185_/A _11185_/B vssd1 vssd1 vccd1 vccd1 _11185_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17801_ _15162_/X _19703_/Q _17805_/S vssd1 vssd1 vccd1 vccd1 _17802_/A sky130_fd_sc_hd__mux2_1
X_10136_ _10175_/A _10135_/X _09621_/X vssd1 vssd1 vccd1 vccd1 _10136_/X sky130_fd_sc_hd__o21a_1
XFILLER_122_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18781_ _19724_/CLK _18781_/D vssd1 vssd1 vccd1 vccd1 _18781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15993_ _15993_/A vssd1 vssd1 vccd1 vccd1 _18995_/D sky130_fd_sc_hd__clkbuf_1
X_17732_ _19681_/Q _17708_/X _17729_/Y _17731_/X vssd1 vssd1 vccd1 vccd1 _19681_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_76_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10067_ _18837_/Q _19391_/Q _19553_/Q _18805_/Q _09808_/A _09936_/A vssd1 vssd1 vccd1
+ vccd1 _10068_/B sky130_fd_sc_hd__mux4_1
X_14944_ _17716_/A _14955_/C vssd1 vssd1 vccd1 vccd1 _14945_/C sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_189_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11122__A3 _18798_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17663_ _17693_/A vssd1 vssd1 vccd1 vccd1 _17686_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_91_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14875_ _14875_/A vssd1 vssd1 vccd1 vccd1 _14875_/X sky130_fd_sc_hd__clkbuf_2
X_19402_ _19660_/CLK _19402_/D vssd1 vssd1 vccd1 vccd1 _19402_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11027__S _11027_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15722__S _15730_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16614_ _16614_/A vssd1 vssd1 vccd1 vccd1 _19262_/D sky130_fd_sc_hd__clkbuf_1
X_13826_ _14102_/A vssd1 vssd1 vccd1 vccd1 _14070_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17594_ _17594_/A vssd1 vssd1 vccd1 vccd1 _19654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19333_ _19397_/CLK _19333_/D vssd1 vssd1 vccd1 vccd1 _19333_/Q sky130_fd_sc_hd__dfxtp_1
X_16545_ _19229_/Q _15548_/X _16547_/S vssd1 vssd1 vccd1 vccd1 _16546_/A sky130_fd_sc_hd__mux2_1
X_13757_ _13686_/X _13606_/X _13757_/S vssd1 vssd1 vccd1 vccd1 _13757_/X sky130_fd_sc_hd__mux2_1
X_10969_ _10969_/A _10969_/B vssd1 vssd1 vccd1 vccd1 _10969_/X sky130_fd_sc_hd__and2_1
X_12708_ _19771_/Q _12666_/B _12707_/X vssd1 vssd1 vccd1 vccd1 _12708_/X sky130_fd_sc_hd__o21a_1
X_19264_ _19818_/CLK _19264_/D vssd1 vssd1 vccd1 vccd1 _19264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11830__A1 _11849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16476_ _16476_/A vssd1 vssd1 vccd1 vccd1 _19198_/D sky130_fd_sc_hd__clkbuf_1
X_13688_ _14192_/B _14093_/A _13689_/S vssd1 vssd1 vccd1 vccd1 _13688_/X sky130_fd_sc_hd__mux2_1
X_18215_ _18223_/A _18215_/B vssd1 vssd1 vccd1 vccd1 _18215_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15427_ _15427_/A vssd1 vssd1 vccd1 vccd1 _18757_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15958__A _17774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12639_ _12639_/A vssd1 vssd1 vccd1 vccd1 _12640_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19195_ _19614_/CLK _19195_/D vssd1 vssd1 vccd1 vccd1 _19195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18146_ _19835_/Q _18148_/C _18145_/Y vssd1 vssd1 vccd1 vccd1 _19835_/D sky130_fd_sc_hd__o21a_1
XFILLER_129_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15358_ _18728_/Q _15162_/X _15362_/S vssd1 vssd1 vccd1 vccd1 _15359_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09882__S0 _09809_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14309_ _14262_/A _14308_/B _13796_/A vssd1 vssd1 vccd1 vccd1 _14309_/X sky130_fd_sc_hd__o21a_1
X_18077_ _18077_/A _18077_/B _18077_/C vssd1 vssd1 vccd1 vccd1 _19812_/D sky130_fd_sc_hd__nor3_1
XANTENNA__16521__A1 _15513_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15289_ _18698_/Q _15168_/X _15289_/S vssd1 vssd1 vccd1 vccd1 _15290_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17028_ _19418_/Q _16689_/X _17036_/S vssd1 vssd1 vccd1 vccd1 _17029_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09850_ _19428_/Q _19204_/Q _19721_/Q _19172_/Q _09914_/A _09843_/A vssd1 vssd1 vccd1
+ vccd1 _09850_/X sky130_fd_sc_hd__mux4_2
XFILLER_124_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09691__A _10417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09781_ _10114_/S vssd1 vssd1 vccd1 vccd1 _09782_/A sky130_fd_sc_hd__clkbuf_4
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ _18982_/CLK _18979_/D vssd1 vssd1 vccd1 vccd1 _18979_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09937__S1 _09936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10321__A1 _11166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15632__S _15636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14063__A2 _14057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12074__A1 _13295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_12_0_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_12_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__11461__A input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09215_ _09215_/A vssd1 vssd1 vccd1 vccd1 _10007_/A sky130_fd_sc_hd__buf_2
XFILLER_167_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09866__A _09866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09146_ _09146_/A vssd1 vssd1 vccd1 vccd1 _09147_/A sky130_fd_sc_hd__buf_4
XFILLER_136_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13388__A _13388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12292__A _19752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16512__A1 _15500_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16699__A _16699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17294__S _17302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10235__S1 _09486_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09979_ _09979_/A vssd1 vssd1 vccd1 vccd1 _09979_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14826__A1 _18436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_190_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _12993_/A _12993_/C _12989_/Y vssd1 vssd1 vccd1 vccd1 _18310_/D sky130_fd_sc_hd__o21a_1
XFILLER_92_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09702__B1 _09184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11941_ _14589_/A _15079_/A vssd1 vssd1 vccd1 vccd1 _11941_/Y sky130_fd_sc_hd__nand2_2
XFILLER_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10312__A1 _19029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _14559_/A _12660_/A _14649_/X input44/X vssd1 vssd1 vccd1 vccd1 _17781_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _11872_/A vssd1 vssd1 vccd1 vccd1 _11879_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__15251__A1 _13149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _13606_/X _13609_/X _13758_/S vssd1 vssd1 vccd1 vccd1 _13611_/X sky130_fd_sc_hd__mux2_1
X_10823_ _10823_/A _10823_/B _10823_/C vssd1 vssd1 vccd1 vccd1 _10823_/X sky130_fd_sc_hd__or3_1
XANTENNA__13570__B _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14591_ _18618_/Q _14591_/B input66/X vssd1 vssd1 vccd1 vccd1 _14680_/A sky130_fd_sc_hd__and3b_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16330_ _16330_/A vssd1 vssd1 vccd1 vccd1 _19134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13542_ _13542_/A _13542_/B vssd1 vssd1 vccd1 vccd1 _13543_/A sky130_fd_sc_hd__and2_1
X_10754_ _19603_/Q _19441_/Q _18887_/Q _18657_/Q _09152_/A _10740_/A vssd1 vssd1 vccd1
+ vccd1 _10755_/B sky130_fd_sc_hd__mux4_1
XFILLER_71_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16261_ _16261_/A vssd1 vssd1 vccd1 vccd1 _19103_/D sky130_fd_sc_hd__clkbuf_1
X_13473_ _18396_/Q _13279_/X _13475_/S vssd1 vssd1 vccd1 vccd1 _13474_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09218__C1 _09217_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10685_ _09179_/A _10684_/X _09209_/A vssd1 vssd1 vccd1 vccd1 _10685_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18000_ _19785_/Q _18000_/B vssd1 vssd1 vccd1 vccd1 _18006_/C sky130_fd_sc_hd__and2_1
X_15212_ _15212_/A vssd1 vssd1 vccd1 vccd1 _18673_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_172_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19638_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12424_ _12424_/A vssd1 vssd1 vccd1 vccd1 _14324_/B sky130_fd_sc_hd__clkbuf_2
X_16192_ _16109_/X _19069_/Q _16194_/S vssd1 vssd1 vccd1 vccd1 _16193_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15143_ _16645_/A vssd1 vssd1 vccd1 vccd1 _15143_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_126_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12355_ _12355_/A vssd1 vssd1 vccd1 vccd1 _14272_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_154_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10474__S1 _09635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11306_ _18425_/Q _18424_/Q vssd1 vssd1 vccd1 vccd1 _11306_/X sky130_fd_sc_hd__or2_1
XFILLER_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12286_ _12286_/A vssd1 vssd1 vccd1 vccd1 _14241_/B sky130_fd_sc_hd__clkbuf_2
X_15074_ _14999_/X _15072_/X _15073_/X vssd1 vssd1 vccd1 vccd1 _16740_/A sky130_fd_sc_hd__o21a_1
XFILLER_107_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_187_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19414_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_141_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15717__S _15719_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18902_ _19295_/CLK _18902_/D vssd1 vssd1 vccd1 vccd1 _18902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14025_ _13975_/X _14024_/Y _13982_/X vssd1 vssd1 vccd1 vccd1 _14025_/Y sky130_fd_sc_hd__a21oi_1
X_11237_ _11239_/A _11235_/C _11235_/A vssd1 vssd1 vccd1 vccd1 _11238_/B sky130_fd_sc_hd__a21oi_1
XFILLER_45_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12930__A _18287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10000__B1 _09231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11168_ _11168_/A _11168_/B vssd1 vssd1 vccd1 vccd1 _11168_/X sky130_fd_sc_hd__or2_1
X_18833_ _19642_/CLK _18833_/D vssd1 vssd1 vccd1 vccd1 _18833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_110_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19082_/CLK sky130_fd_sc_hd__clkbuf_16
X_10119_ _18772_/Q _19001_/Q _18932_/Q _19230_/Q _10011_/S _09147_/A vssd1 vssd1 vccd1
+ vccd1 _10120_/B sky130_fd_sc_hd__mux4_1
XFILLER_96_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18764_ _19707_/CLK _18764_/D vssd1 vssd1 vccd1 vccd1 _18764_/Q sky130_fd_sc_hd__dfxtp_1
X_15976_ _15976_/A vssd1 vssd1 vccd1 vccd1 _18987_/D sky130_fd_sc_hd__clkbuf_1
X_11099_ _11099_/A _11099_/B vssd1 vssd1 vccd1 vccd1 _11099_/X sky130_fd_sc_hd__or2_1
X_17715_ _19678_/Q _17708_/X _17712_/Y _17714_/X vssd1 vssd1 vccd1 vccd1 _19678_/D
+ sky130_fd_sc_hd__o22a_1
X_14927_ _11542_/X _14923_/X _14926_/X vssd1 vssd1 vccd1 vccd1 _16699_/A sky130_fd_sc_hd__o21a_2
X_18695_ _19571_/CLK _18695_/D vssd1 vssd1 vccd1 vccd1 _18695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13761__A _13761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17646_ _13230_/X _17645_/Y _17658_/S vssd1 vssd1 vccd1 vccd1 _17646_/X sky130_fd_sc_hd__mux2_1
X_14858_ _14858_/A vssd1 vssd1 vccd1 vccd1 _18598_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_125_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19686_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09450__S _10348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13809_ _13891_/A vssd1 vssd1 vccd1 vccd1 _13810_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17577_ _19647_/Q _16803_/A _17579_/S vssd1 vssd1 vccd1 vccd1 _17578_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14789_ _14787_/Y _14788_/X _14893_/A vssd1 vssd1 vccd1 vccd1 _14789_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19316_ _19639_/CLK _19316_/D vssd1 vssd1 vccd1 vccd1 _19316_/Q sky130_fd_sc_hd__dfxtp_1
X_16528_ _19221_/Q _15522_/X _16536_/S vssd1 vssd1 vccd1 vccd1 _16529_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12096__B _12096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10162__S0 _10200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17379__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15688__A _15734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19247_ _19633_/CLK _19247_/D vssd1 vssd1 vccd1 vccd1 _19247_/Q sky130_fd_sc_hd__dfxtp_1
X_16459_ _16459_/A vssd1 vssd1 vccd1 vccd1 _19190_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16283__S _16283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13556__A1 _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19178_ _19660_/CLK _19178_/D vssd1 vssd1 vccd1 vccd1 _19178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09855__S0 _09163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18129_ _18173_/A vssd1 vssd1 vccd1 vccd1 _18165_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_117_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09902_ _19524_/Q _19138_/Q _19588_/Q _18744_/Q _09782_/X _09783_/X vssd1 vssd1 vccd1
+ vccd1 _09903_/B sky130_fd_sc_hd__mux4_2
XFILLER_132_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09833_ _10044_/A vssd1 vssd1 vccd1 vccd1 _09879_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09764_ _19267_/Q _19038_/Q _18969_/Q _19363_/Q _09760_/X _09763_/X vssd1 vssd1 vccd1
+ vccd1 _09764_/X sky130_fd_sc_hd__mux4_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12295__A1 _19683_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16458__S _16464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09695_ _09695_/A vssd1 vssd1 vccd1 vccd1 _09704_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13671__A _13671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15362__S _15362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12047__A1 _19673_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14992__A0 _18450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11622__C _13671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17289__S _17291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_137_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09596__A _10400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10470_ _18764_/Q _18993_/Q _18924_/Q _19222_/Q _10560_/S _09634_/A vssd1 vssd1 vccd1
+ vccd1 _10471_/B sky130_fd_sc_hd__mux4_1
XFILLER_136_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09129_ _19695_/Q vssd1 vssd1 vccd1 vccd1 _10823_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12140_ _12089_/A _12089_/B _12114_/A _12139_/X vssd1 vssd1 vccd1 vccd1 _12141_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_155_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10781__A1 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12071_ _19674_/Q _12412_/B vssd1 vssd1 vccd1 vccd1 _12071_/X sky130_fd_sc_hd__or2_1
XFILLER_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11022_ _18427_/Q vssd1 vssd1 vccd1 vccd1 _11022_/X sky130_fd_sc_hd__buf_6
XFILLER_104_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15830_ _14821_/X _18922_/Q _15830_/S vssd1 vssd1 vccd1 vccd1 _15831_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17749__A0 _19685_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15761_ _14833_/X _18891_/Q _15769_/S vssd1 vssd1 vccd1 vccd1 _15762_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12973_ _12983_/A _12973_/B _12973_/C vssd1 vssd1 vccd1 vccd1 _18305_/D sky130_fd_sc_hd__nor3_1
XFILLER_18_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_42_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19657_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14677__A _14677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15272__S _15278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17500_ _17500_/A vssd1 vssd1 vccd1 vccd1 _19612_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ input1/X _14703_/X _14708_/X _14711_/X vssd1 vssd1 vccd1 vccd1 _16639_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10297__B1 _09625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _11879_/A _11879_/B _11899_/A _11923_/Y vssd1 vssd1 vccd1 vccd1 _11925_/B
+ sky130_fd_sc_hd__a31o_2
X_18480_ _18482_/CLK _18480_/D vssd1 vssd1 vccd1 vccd1 _18480_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _15692_/A vssd1 vssd1 vccd1 vccd1 _18860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17431_ _16800_/X _19582_/Q _17435_/S vssd1 vssd1 vccd1 vccd1 _17432_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _18205_/A vssd1 vssd1 vccd1 vccd1 _14643_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11855_ _18356_/Q _11820_/B _11825_/X vssd1 vssd1 vccd1 vccd1 _11888_/D sky130_fd_sc_hd__a21bo_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output105_A _09106_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10806_ _19601_/Q _19439_/Q _18885_/Q _18655_/Q _10932_/S _10713_/A vssd1 vssd1 vccd1
+ vccd1 _10807_/B sky130_fd_sc_hd__mux4_1
XFILLER_32_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17362_ _17362_/A vssd1 vssd1 vccd1 vccd1 _19551_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_57_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19329_/CLK sky130_fd_sc_hd__clkbuf_16
X_14574_ _18546_/Q _14564_/X _14572_/Y _14573_/X vssd1 vssd1 vccd1 vccd1 _18546_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18174__B1 _19845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11786_ _11785_/Y _11747_/B _11745_/A vssd1 vssd1 vccd1 vccd1 _11787_/B sky130_fd_sc_hd__o21a_2
X_19101_ _19647_/CLK _19101_/D vssd1 vssd1 vccd1 vccd1 _19101_/Q sky130_fd_sc_hd__dfxtp_1
X_16313_ _16313_/A vssd1 vssd1 vccd1 vccd1 _19126_/D sky130_fd_sc_hd__clkbuf_1
X_13525_ _13525_/A _14431_/C vssd1 vssd1 vccd1 vccd1 _13545_/C sky130_fd_sc_hd__nor2_1
X_17293_ _17304_/A vssd1 vssd1 vccd1 vccd1 _17302_/S sky130_fd_sc_hd__clkbuf_8
X_10737_ _10982_/S vssd1 vssd1 vccd1 vccd1 _10858_/A sky130_fd_sc_hd__buf_2
XFILLER_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19032_ _19647_/CLK _19032_/D vssd1 vssd1 vccd1 vccd1 _19032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16244_ _16077_/X _19096_/Q _16246_/S vssd1 vssd1 vccd1 vccd1 _16245_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13538__B2 _12555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13456_ _18388_/Q _13197_/X _13464_/S vssd1 vssd1 vccd1 vccd1 _13457_/A sky130_fd_sc_hd__mux2_1
X_10668_ _10668_/A vssd1 vssd1 vccd1 vccd1 _10669_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12407_ _12408_/B vssd1 vssd1 vccd1 vccd1 _12407_/Y sky130_fd_sc_hd__inv_2
X_16175_ _16083_/X _19061_/Q _16183_/S vssd1 vssd1 vccd1 vccd1 _16176_/A sky130_fd_sc_hd__mux2_1
X_13387_ _12577_/X _13379_/Y _13386_/X _12596_/X _18646_/Q vssd1 vssd1 vccd1 vccd1
+ _13387_/X sky130_fd_sc_hd__a32o_4
XFILLER_12_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10599_ _09927_/A _10589_/X _10598_/X _09307_/A _18435_/Q vssd1 vssd1 vccd1 vccd1
+ _12474_/B sky130_fd_sc_hd__a32o_4
XANTENNA__10221__A0 _19614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput107 _13570_/B vssd1 vssd1 vccd1 vccd1 io_dbus_ld_type[2] sky130_fd_sc_hd__buf_2
XFILLER_114_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15126_ _18644_/Q _15123_/X _15125_/X _09898_/A vssd1 vssd1 vccd1 vccd1 _18644_/D
+ sky130_fd_sc_hd__a22o_1
Xoutput118 _12485_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[16] sky130_fd_sc_hd__buf_2
XFILLER_142_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12338_ _19685_/Q _13529_/B vssd1 vssd1 vccd1 vccd1 _12338_/X sky130_fd_sc_hd__or2_1
Xoutput129 _12500_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[26] sky130_fd_sc_hd__buf_2
XFILLER_142_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15057_ _15057_/A vssd1 vssd1 vccd1 vccd1 _18615_/D sky130_fd_sc_hd__clkbuf_1
X_12269_ _12265_/Y _12268_/Y _12389_/S vssd1 vssd1 vccd1 vccd1 _12269_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12660__A _12660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14008_ _14005_/B _13658_/X _14276_/A vssd1 vssd1 vccd1 vccd1 _14008_/X sky130_fd_sc_hd__a21o_1
X_19865_ _19866_/CLK _19865_/D vssd1 vssd1 vccd1 vccd1 _19865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18816_ _19648_/CLK _18816_/D vssd1 vssd1 vccd1 vccd1 _18816_/Q sky130_fd_sc_hd__dfxtp_1
X_19796_ _19798_/CLK _19796_/D vssd1 vssd1 vccd1 vccd1 _19796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18747_ _19722_/CLK _18747_/D vssd1 vssd1 vccd1 vccd1 _18747_/Q sky130_fd_sc_hd__dfxtp_1
X_15959_ _17774_/A _15959_/B vssd1 vssd1 vccd1 vccd1 _18981_/D sky130_fd_sc_hd__nor2_2
XANTENNA__14587__A _14587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15182__S _15185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09480_ _09480_/A vssd1 vssd1 vccd1 vccd1 _09481_/A sky130_fd_sc_hd__buf_4
X_18678_ _19592_/CLK _18678_/D vssd1 vssd1 vccd1 vccd1 _18678_/Q sky130_fd_sc_hd__dfxtp_1
X_17629_ _17707_/A vssd1 vssd1 vccd1 vccd1 _17653_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_36_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10135__S0 _09729_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10686__S1 _09139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12554__B _12554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12201__A1 _19748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16741__S _16741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__A _11088_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16977__A _16977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09816_ _09819_/A _09815_/X _09320_/X vssd1 vssd1 vccd1 vccd1 _09816_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_100_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_63_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09747_ _10144_/A _09747_/B vssd1 vssd1 vccd1 vccd1 _09747_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16188__S _16194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09678_ _18780_/Q _19009_/Q _18940_/Q _19238_/Q _09600_/A _10280_/A vssd1 vssd1 vccd1
+ vccd1 _09678_/X sky130_fd_sc_hd__mux4_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10374__S0 _09448_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11640_/A _11640_/B vssd1 vssd1 vccd1 vccd1 _11640_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11571_ _19728_/Q _17855_/C vssd1 vssd1 vccd1 vccd1 _11572_/A sky130_fd_sc_hd__and2_1
XFILLER_156_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13310_ _13267_/X _13307_/X _13309_/X _13282_/X vssd1 vssd1 vccd1 vccd1 _18365_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_168_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10522_ _09679_/A _10521_/X _10219_/A vssd1 vssd1 vccd1 vccd1 _10522_/X sky130_fd_sc_hd__o21a_1
XFILLER_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14290_ _13806_/X _14288_/B _14289_/X _14000_/X vssd1 vssd1 vccd1 vccd1 _14290_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13241_ _19865_/Q _12525_/X _12736_/A _19833_/Q vssd1 vssd1 vccd1 vccd1 _14813_/C
+ sky130_fd_sc_hd__a22o_2
XFILLER_155_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10453_ _18765_/Q _18994_/Q _18925_/Q _19223_/Q _10224_/X _11111_/A vssd1 vssd1 vccd1
+ vccd1 _10453_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13172_ _18271_/Q _13404_/B vssd1 vssd1 vccd1 vccd1 _13172_/X sky130_fd_sc_hd__and2_1
XFILLER_164_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input66_A io_ibus_valid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ _10384_/A vssd1 vssd1 vccd1 vccd1 _10384_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12123_ _18367_/Q _18366_/Q _12123_/C vssd1 vssd1 vccd1 vccd1 _12169_/C sky130_fd_sc_hd__and3_1
X_17980_ _17980_/A _17980_/B _17981_/B vssd1 vssd1 vccd1 vccd1 _19778_/D sky130_fd_sc_hd__nor3_1
XFILLER_151_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12480__A _12480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16931_ _16758_/X _19375_/Q _16931_/S vssd1 vssd1 vccd1 vccd1 _16932_/A sky130_fd_sc_hd__mux2_1
X_12054_ _11497_/A _12026_/X _12126_/A _12483_/A vssd1 vssd1 vccd1 vccd1 _12055_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10506__A1 _09927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10506__B2 _18437_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11005_ _10772_/A _11004_/X _11065_/A vssd1 vssd1 vccd1 vccd1 _11005_/X sky130_fd_sc_hd__a21o_1
XFILLER_78_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19650_ _19812_/CLK _19650_/D vssd1 vssd1 vccd1 vccd1 _19650_/Q sky130_fd_sc_hd__dfxtp_1
X_16862_ _16862_/A vssd1 vssd1 vccd1 vccd1 _19344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15813_ _14729_/X _18914_/Q _15819_/S vssd1 vssd1 vccd1 vccd1 _15814_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18601_ _19580_/CLK _18601_/D vssd1 vssd1 vccd1 vccd1 _18601_/Q sky130_fd_sc_hd__dfxtp_1
X_19581_ _19581_/CLK _19581_/D vssd1 vssd1 vccd1 vccd1 _19581_/Q sky130_fd_sc_hd__dfxtp_1
X_16793_ _16793_/A vssd1 vssd1 vccd1 vccd1 _16793_/X sky130_fd_sc_hd__clkbuf_2
X_18532_ _18618_/CLK _18532_/D vssd1 vssd1 vccd1 vccd1 _18532_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15744_ _15744_/A vssd1 vssd1 vccd1 vccd1 _18883_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12956_ _18295_/Q _12957_/C _18296_/Q vssd1 vssd1 vccd1 vccd1 _12958_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__17198__A1 _12598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ _13246_/A _11962_/D vssd1 vssd1 vccd1 vccd1 _11907_/X sky130_fd_sc_hd__or2_1
X_18463_ _19693_/CLK _18463_/D vssd1 vssd1 vccd1 vccd1 _18463_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15675_ _18853_/Q _15503_/X _15675_/S vssd1 vssd1 vccd1 vccd1 _15676_/A sky130_fd_sc_hd__mux2_1
X_12887_ _12897_/A _12893_/C vssd1 vssd1 vccd1 vccd1 _12887_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17414_ _17414_/A vssd1 vssd1 vccd1 vccd1 _19574_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15730__S _15730_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _14696_/A vssd1 vssd1 vccd1 vccd1 _14654_/A sky130_fd_sc_hd__buf_2
XFILLER_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11219__C1 _11204_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18394_ _18395_/CLK _18394_/D vssd1 vssd1 vccd1 vccd1 _18394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11838_ _11940_/A _11939_/B vssd1 vssd1 vccd1 vccd1 _11839_/B sky130_fd_sc_hd__nand2_2
XANTENNA__14956__B1 _14744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17345_ _17345_/A vssd1 vssd1 vccd1 vccd1 _19543_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _14557_/A _14559_/B vssd1 vssd1 vccd1 vccd1 _14557_/X sky130_fd_sc_hd__or2_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11769_ _11768_/A _11768_/B _11827_/B vssd1 vssd1 vccd1 vccd1 _11769_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13508_ _18412_/Q _13412_/X _13508_/S vssd1 vssd1 vccd1 vccd1 _13509_/A sky130_fd_sc_hd__mux2_1
X_17276_ _19513_/Q _16680_/X _17280_/S vssd1 vssd1 vccd1 vccd1 _17277_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14488_ _14488_/A vssd1 vssd1 vccd1 vccd1 _18514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19015_ _19632_/CLK _19015_/D vssd1 vssd1 vccd1 vccd1 _19015_/Q sky130_fd_sc_hd__dfxtp_1
X_16227_ _16051_/X _19088_/Q _16235_/S vssd1 vssd1 vccd1 vccd1 _16228_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13439_ _13311_/A _13437_/Y _13438_/X _13401_/X vssd1 vssd1 vccd1 vccd1 _18381_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16561__S _16569_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16158_ _16158_/A vssd1 vssd1 vccd1 vccd1 _19053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15109_ _15116_/A vssd1 vssd1 vccd1 vccd1 _15109_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12390__A _19687_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16089_ _16089_/A vssd1 vssd1 vccd1 vccd1 _19030_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10903__A _18428_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10840__S1 _10713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15684__A1 _15516_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15905__S _15913_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19848_ _19851_/CLK _19848_/D vssd1 vssd1 vccd1 vccd1 _19848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09601_ _10384_/A vssd1 vssd1 vccd1 vccd1 _09602_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19779_ _19779_/CLK _19779_/D vssd1 vssd1 vccd1 vccd1 _19779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09532_ _09519_/X _09531_/X _10494_/A vssd1 vssd1 vccd1 vccd1 _09532_/X sky130_fd_sc_hd__mux2_2
XFILLER_71_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11453__B _14431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ _09463_/A _09463_/B vssd1 vssd1 vccd1 vccd1 _09463_/X sky130_fd_sc_hd__or2_1
XFILLER_25_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09394_ _09394_/A vssd1 vssd1 vccd1 vccd1 _09395_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17897__C1 _14585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14175__A1 _18443_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14175__B2 _14174_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10085__A _10262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12725__A2 _12665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11933__B1 _14431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10831__S1 _10740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10813__A _10813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15675__A1 _15503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13686__A0 _14155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15815__S _15819_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12810_ _12810_/A vssd1 vssd1 vccd1 vccd1 _18034_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13989__A1 _11813_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15116__A _15116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13790_ _13879_/S vssd1 vssd1 vccd1 vccd1 _13880_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__09657__A2 _09647_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _13235_/A vssd1 vssd1 vccd1 vccd1 _12741_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10898__S1 _10785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _15460_/A vssd1 vssd1 vccd1 vccd1 _18772_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _19472_/Q _13235_/A _12671_/X _18687_/Q vssd1 vssd1 vccd1 vccd1 _12672_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _14411_/A vssd1 vssd1 vccd1 vccd1 _18482_/D sky130_fd_sc_hd__clkbuf_1
X_11623_ _11621_/X _11623_/B vssd1 vssd1 vccd1 vccd1 _11624_/B sky130_fd_sc_hd__and2b_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15391_ _18743_/Q _15210_/X _15395_/S vssd1 vssd1 vccd1 vccd1 _15392_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17130_ _16838_/X _19464_/Q _17130_/S vssd1 vssd1 vccd1 vccd1 _17131_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14342_ _14342_/A vssd1 vssd1 vccd1 vccd1 _18458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11554_ _11554_/A vssd1 vssd1 vccd1 vccd1 _19081_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10505_ _09412_/A _10496_/X _10498_/X _10504_/X _09392_/A vssd1 vssd1 vccd1 vccd1
+ _10505_/X sky130_fd_sc_hd__a311o_4
X_17061_ _17061_/A vssd1 vssd1 vccd1 vccd1 _19433_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17477__S _17485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14273_ _13977_/A _14272_/B _14040_/A vssd1 vssd1 vccd1 vccd1 _14273_/X sky130_fd_sc_hd__o21a_1
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11485_ _11485_/A vssd1 vssd1 vccd1 vccd1 _11550_/B sky130_fd_sc_hd__buf_2
XFILLER_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16012_ _14975_/X _19004_/Q _16016_/S vssd1 vssd1 vccd1 vccd1 _16013_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13224_ _18358_/Q _13127_/A _13221_/X _13223_/X vssd1 vssd1 vccd1 vccd1 _13224_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12716__A2 _12713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10436_ _09275_/A _10426_/X _10435_/X _09282_/A _18438_/Q vssd1 vssd1 vccd1 vccd1
+ _10461_/A sky130_fd_sc_hd__a32o_4
XFILLER_152_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13155_ _19471_/Q _13235_/A _12671_/X _18686_/Q vssd1 vssd1 vccd1 vccd1 _13155_/X
+ sky130_fd_sc_hd__a22o_1
X_10367_ _10367_/A vssd1 vssd1 vccd1 vccd1 _10368_/A sky130_fd_sc_hd__buf_4
XANTENNA__10723__A _10797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _12106_/A vssd1 vssd1 vccd1 vccd1 _13567_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17963_ _19772_/Q _19771_/Q _17963_/C vssd1 vssd1 vccd1 vccd1 _17965_/B sky130_fd_sc_hd__and3_1
X_13086_ _18626_/Q _13086_/B vssd1 vssd1 vccd1 vccd1 _13086_/X sky130_fd_sc_hd__or2_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _10299_/A _12485_/A vssd1 vssd1 vccd1 vccd1 _10300_/A sky130_fd_sc_hd__and2_1
XANTENNA__13141__A2 _13235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19702_ _19702_/CLK _19702_/D vssd1 vssd1 vccd1 vccd1 _19702_/Q sky130_fd_sc_hd__dfxtp_1
X_12037_ _11975_/A _12011_/A _12010_/A _13595_/A vssd1 vssd1 vccd1 vccd1 _12037_/X
+ sky130_fd_sc_hd__a22o_1
X_16914_ _16914_/A vssd1 vssd1 vccd1 vccd1 _19368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17894_ _17894_/A vssd1 vssd1 vccd1 vccd1 _19747_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15418__A1 _15133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10586__S0 _10500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19633_ _19633_/CLK _19633_/D vssd1 vssd1 vccd1 vccd1 _19633_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13429__B1 _12671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16845_ _16844_/X _19338_/Q _16845_/S vssd1 vssd1 vccd1 vccd1 _16846_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19564_ _19648_/CLK _19564_/D vssd1 vssd1 vccd1 vccd1 _19564_/Q sky130_fd_sc_hd__dfxtp_1
X_16776_ _16776_/A vssd1 vssd1 vccd1 vccd1 _19316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13988_ _13738_/X _13970_/X _13987_/X _13784_/X vssd1 vssd1 vccd1 vccd1 _13988_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10338__S0 _11188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18515_ _18519_/CLK _18515_/D vssd1 vssd1 vccd1 vccd1 _18515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15727_ _15727_/A vssd1 vssd1 vccd1 vccd1 _18876_/D sky130_fd_sc_hd__clkbuf_1
X_12939_ _18290_/Q _18289_/Q _12939_/C vssd1 vssd1 vccd1 vccd1 _12946_/C sky130_fd_sc_hd__and3_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16556__S _16558_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19495_ _19795_/CLK _19495_/D vssd1 vssd1 vccd1 vccd1 _19495_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10112__C1 _09249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10889__S1 _10785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18446_ _19695_/CLK _18446_/D vssd1 vssd1 vccd1 vccd1 _18446_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_61_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15658_ _18846_/Q _15583_/X _15658_/S vssd1 vssd1 vccd1 vccd1 _15659_/A sky130_fd_sc_hd__mux2_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14609_ _14609_/A vssd1 vssd1 vccd1 vccd1 _18557_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18377_ _19690_/CLK _18377_/D vssd1 vssd1 vccd1 vccd1 _18377_/Q sky130_fd_sc_hd__dfxtp_1
X_15589_ _16844_/A vssd1 vssd1 vccd1 vccd1 _15589_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17328_ _16755_/X _19536_/Q _17330_/S vssd1 vssd1 vccd1 vccd1 _17329_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17879__C1 _12802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17387__S _17389_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17259_ _17259_/A vssd1 vssd1 vccd1 vccd1 _19505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09694__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10633__A _10785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13668__A0 _12381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09515_ _09515_/A vssd1 vssd1 vccd1 vccd1 _09587_/A sky130_fd_sc_hd__clkbuf_4
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09869__A _09869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _09449_/A vssd1 vssd1 vccd1 vccd1 _09447_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09377_ _10762_/A vssd1 vssd1 vccd1 vccd1 _10593_/A sky130_fd_sc_hd__buf_2
XFILLER_40_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14148__A1 _12066_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11270_ _11269_/B _11269_/C _11269_/A vssd1 vssd1 vccd1 vccd1 _11271_/B sky130_fd_sc_hd__a21o_1
XFILLER_118_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10221_ _19614_/Q _19452_/Q _18898_/Q _18668_/Q _09673_/S _09602_/A vssd1 vssd1 vccd1
+ vccd1 _10222_/B sky130_fd_sc_hd__mux4_1
XFILLER_161_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10804__S1 _10726_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11382__B2 _18417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ _10167_/A _10152_/B vssd1 vssd1 vccd1 vccd1 _10152_/X sky130_fd_sc_hd__or2_1
XANTENNA__13659__A0 _12282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10083_ _10093_/A _10079_/X _10082_/X _09230_/A vssd1 vssd1 vccd1 vccd1 _10083_/X
+ sky130_fd_sc_hd__o211a_1
X_14960_ _14960_/A vssd1 vssd1 vccd1 vccd1 _14960_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09422__S1 _09364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13911_ _11704_/Y _13827_/X _13828_/X vssd1 vssd1 vccd1 vccd1 _13911_/X sky130_fd_sc_hd__a21o_1
XFILLER_47_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input29_A io_dbus_rdata[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14891_ _14889_/X _18601_/Q _14941_/S vssd1 vssd1 vccd1 vccd1 _14892_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16630_ _16630_/A vssd1 vssd1 vccd1 vccd1 _19270_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13842_ _14135_/A _13841_/X _13810_/A vssd1 vssd1 vccd1 vccd1 _13842_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16561_ _19236_/Q _15570_/X _16569_/S vssd1 vssd1 vccd1 vccd1 _16562_/A sky130_fd_sc_hd__mux2_1
X_13773_ _13771_/X _13772_/X _13776_/S vssd1 vssd1 vccd1 vccd1 _13773_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10985_ _10548_/A _10982_/X _10984_/X vssd1 vssd1 vccd1 vccd1 _10985_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18300_ _19856_/CLK _18300_/D vssd1 vssd1 vccd1 vccd1 _18300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15512_ _15512_/A vssd1 vssd1 vccd1 vccd1 _18791_/D sky130_fd_sc_hd__clkbuf_1
X_12724_ _19868_/Q _12604_/X _12528_/A _19836_/Q _12723_/X vssd1 vssd1 vccd1 vccd1
+ _12724_/X sky130_fd_sc_hd__a221o_2
X_19280_ _19506_/CLK _19280_/D vssd1 vssd1 vccd1 vccd1 _19280_/Q sky130_fd_sc_hd__dfxtp_1
X_16492_ _16492_/A vssd1 vssd1 vccd1 vccd1 _19205_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18231_ _19865_/Q _19864_/Q _18231_/C vssd1 vssd1 vccd1 vccd1 _18232_/B sky130_fd_sc_hd__and3_1
X_15443_ _15443_/A vssd1 vssd1 vccd1 vccd1 _18764_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12655_ _12600_/X _12636_/Y _12654_/X _12558_/X _18639_/Q vssd1 vssd1 vccd1 vccd1
+ _12656_/B sky130_fd_sc_hd__a32o_4
XFILLER_169_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10718__A _10807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18162_ _19841_/Q _18164_/C _18161_/Y vssd1 vssd1 vccd1 vccd1 _19841_/D sky130_fd_sc_hd__o21a_1
X_11606_ _11357_/Y _11584_/A _11644_/B _13570_/D _13585_/B vssd1 vssd1 vccd1 vccd1
+ _11606_/X sky130_fd_sc_hd__a2111o_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15374_ _15374_/A vssd1 vssd1 vccd1 vccd1 _18735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12586_ _18284_/Q _12606_/A _12642_/A _18367_/Q vssd1 vssd1 vccd1 vccd1 _12586_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10948__A1 _10950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17113_ _16813_/X _19456_/Q _17119_/S vssd1 vssd1 vccd1 vccd1 _17114_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_185_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14325_ _13806_/X _14323_/B _14324_/X _14000_/X vssd1 vssd1 vccd1 vccd1 _14325_/X
+ sky130_fd_sc_hd__o211a_1
X_18093_ _18094_/A _18094_/C _18092_/Y vssd1 vssd1 vccd1 vccd1 _19817_/D sky130_fd_sc_hd__o21a_1
XFILLER_128_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11537_ _13570_/A _11360_/C _12277_/B _11537_/D vssd1 vssd1 vccd1 vccd1 _11538_/D
+ sky130_fd_sc_hd__and4bb_1
XFILLER_172_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12933__A _18288_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17044_ _17044_/A vssd1 vssd1 vccd1 vccd1 _19425_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_output97_A _12450_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14256_ _14037_/X _13999_/X _14255_/Y _13737_/A vssd1 vssd1 vccd1 vccd1 _14256_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11468_ _14524_/A _11468_/B _11468_/C vssd1 vssd1 vccd1 vccd1 _11966_/B sky130_fd_sc_hd__and3_2
X_13207_ _19798_/Q _12748_/A _12752_/A _19766_/Q vssd1 vssd1 vccd1 vccd1 _13207_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10419_ _09171_/A _10418_/X _11099_/A vssd1 vssd1 vccd1 vccd1 _10419_/X sky130_fd_sc_hd__a21o_1
XFILLER_48_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14187_ _14187_/A vssd1 vssd1 vccd1 vccd1 _18444_/D sky130_fd_sc_hd__clkbuf_1
X_11399_ _11400_/A _11404_/A _11401_/A vssd1 vssd1 vccd1 vccd1 _12639_/A sky130_fd_sc_hd__nor3_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _18350_/Q _13118_/X _13137_/X vssd1 vssd1 vccd1 vccd1 _18350_/D sky130_fd_sc_hd__a21o_1
XFILLER_98_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18977__D _18977_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18995_ _19707_/CLK _18995_/D vssd1 vssd1 vccd1 vccd1 _18995_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15455__S _15459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17946_ _19767_/Q _19766_/Q _19765_/Q _17946_/D vssd1 vssd1 vccd1 vccd1 _17957_/D
+ sky130_fd_sc_hd__and4_1
X_13069_ _18332_/Q _18331_/Q _18333_/Q _13069_/D vssd1 vssd1 vccd1 vccd1 _18112_/D
+ sky130_fd_sc_hd__and4_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12322__B1 _19753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17877_ _17877_/A vssd1 vssd1 vccd1 vccd1 _19739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19616_ _19616_/CLK _19616_/D vssd1 vssd1 vccd1 vccd1 _19616_/Q sky130_fd_sc_hd__dfxtp_1
X_16828_ _16828_/A vssd1 vssd1 vccd1 vccd1 _19332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19547_ _19579_/CLK _19547_/D vssd1 vssd1 vccd1 vccd1 _19547_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12625__B2 _19488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16759_ _16758_/X _19311_/Q _16759_/S vssd1 vssd1 vccd1 vccd1 _16760_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09300_ _18577_/Q vssd1 vssd1 vccd1 vccd1 _13523_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09689__A _09689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19478_ _19488_/CLK _19478_/D vssd1 vssd1 vccd1 vccd1 _19478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17564__A1 _16784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09231_ _09231_/A vssd1 vssd1 vccd1 vccd1 _09231_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__14378__A1 _18503_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18429_ _18982_/CLK _18429_/D vssd1 vssd1 vccd1 vccd1 _18429_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12389__A0 _12385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13004__A _13034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09162_ _09911_/S vssd1 vssd1 vccd1 vccd1 _09163_/A sky130_fd_sc_hd__buf_4
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10347__B _12483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09093_ _13526_/A _12471_/B _11313_/D vssd1 vssd1 vccd1 vccd1 _09094_/A sky130_fd_sc_hd__nor3_4
XFILLER_163_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12562__B _13042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16034__B _17064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13353__A2 _13139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17845__S _17849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09995_ _09995_/A vssd1 vssd1 vccd1 vccd1 _09996_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_131_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15365__S _15373_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13105__A2 _12731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11116__A1 _10447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09599__A _10279_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ _18592_/Q _19281_/Q _10770_/S vssd1 vssd1 vccd1 vccd1 _10770_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09429_ _09429_/A vssd1 vssd1 vccd1 vccd1 _09430_/A sky130_fd_sc_hd__buf_2
XFILLER_139_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12440_ _12196_/X _12438_/X _12455_/B _11801_/X vssd1 vssd1 vccd1 vccd1 _12440_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_139_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12371_ _12371_/A _12371_/B _12371_/C vssd1 vssd1 vccd1 vccd1 _12371_/X sky130_fd_sc_hd__and3_1
XFILLER_139_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14110_ _14088_/X _14107_/X _14109_/X vssd1 vssd1 vccd1 vccd1 _14110_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09891__S1 _09881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11322_ _11337_/A _14524_/A _11343_/C _11322_/D vssd1 vssd1 vccd1 vccd1 _11372_/B
+ sky130_fd_sc_hd__and4_1
X_15090_ _18622_/Q _15089_/X _15093_/S vssd1 vssd1 vccd1 vccd1 _15091_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09548__A1 _09978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14041_ _14059_/A _14045_/A _14040_/X vssd1 vssd1 vccd1 vccd1 _14041_/X sky130_fd_sc_hd__o21a_1
X_11253_ _11047_/X _12458_/A _11024_/X vssd1 vssd1 vccd1 vccd1 _11253_/X sky130_fd_sc_hd__o21a_1
XFILLER_107_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10204_ _19420_/Q _19196_/Q _19713_/Q _19164_/Q _09795_/A _10080_/X vssd1 vssd1 vccd1
+ vccd1 _10204_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11184_ _19271_/Q _19042_/Q _18973_/Q _19367_/Q _10129_/S _09736_/A vssd1 vssd1 vccd1
+ vccd1 _11185_/B sky130_fd_sc_hd__mux4_1
X_17800_ _17800_/A vssd1 vssd1 vccd1 vccd1 _19702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10135_ _19422_/Q _19198_/Q _19715_/Q _19166_/Q _09729_/S _10331_/A vssd1 vssd1 vccd1
+ vccd1 _10135_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15992_ _14867_/X _18995_/Q _15994_/S vssd1 vssd1 vccd1 vccd1 _15993_/A sky130_fd_sc_hd__mux2_1
X_18780_ _19723_/CLK _18780_/D vssd1 vssd1 vccd1 vccd1 _18780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10066_ _10044_/A _10065_/X _09892_/A vssd1 vssd1 vccd1 vccd1 _10066_/X sky130_fd_sc_hd__o21a_1
X_17731_ _17730_/X _13346_/X _17724_/X vssd1 vssd1 vccd1 vccd1 _17731_/X sky130_fd_sc_hd__a21bo_1
X_14943_ _17716_/A _14955_/C vssd1 vssd1 vccd1 vccd1 _14943_/X sky130_fd_sc_hd__and2_1
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17490__S _17496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09720__B2 _18452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17662_ _17662_/A _17667_/C vssd1 vssd1 vccd1 vccd1 _17662_/Y sky130_fd_sc_hd__xnor2_2
X_14874_ _18440_/Q _14839_/S _14873_/X vssd1 vssd1 vccd1 vccd1 _14874_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10961__S0 _10959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19401_ _19595_/CLK _19401_/D vssd1 vssd1 vccd1 vccd1 _19401_/Q sky130_fd_sc_hd__dfxtp_1
X_16613_ _19262_/Q vssd1 vssd1 vccd1 vccd1 _16614_/A sky130_fd_sc_hd__clkbuf_1
X_13825_ _13738_/X _13782_/X _13784_/X _13824_/X vssd1 vssd1 vccd1 vccd1 _13825_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17593_ _19654_/Q _16825_/A _17601_/S vssd1 vssd1 vccd1 vccd1 _17594_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19332_ _19622_/CLK _19332_/D vssd1 vssd1 vccd1 vccd1 _19332_/Q sky130_fd_sc_hd__dfxtp_1
X_16544_ _16544_/A vssd1 vssd1 vccd1 vccd1 _19228_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13756_ _13754_/X _13755_/X _13759_/S vssd1 vssd1 vccd1 vccd1 _13756_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10968_ _18589_/Q _19278_/Q _10983_/S vssd1 vssd1 vccd1 vccd1 _10969_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12707_ _19670_/Q _12737_/A _12706_/X vssd1 vssd1 vccd1 vccd1 _12707_/X sky130_fd_sc_hd__a21o_1
X_19263_ _19810_/CLK _19263_/D vssd1 vssd1 vccd1 vccd1 _19263_/Q sky130_fd_sc_hd__dfxtp_1
X_16475_ _16096_/X _19198_/Q _16475_/S vssd1 vssd1 vccd1 vccd1 _16476_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13687_ _13685_/X _13686_/X _13757_/S vssd1 vssd1 vccd1 vccd1 _13687_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10899_ _10899_/A _10899_/B vssd1 vssd1 vccd1 vccd1 _10899_/Y sky130_fd_sc_hd__nor2_1
X_18214_ _19859_/Q _18214_/B _18214_/C vssd1 vssd1 vccd1 vccd1 _18215_/B sky130_fd_sc_hd__and3_1
X_15426_ _18757_/Q _15152_/X _15426_/S vssd1 vssd1 vccd1 vccd1 _15427_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12638_ _13270_/B vssd1 vssd1 vccd1 vccd1 _12638_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19194_ _19647_/CLK _19194_/D vssd1 vssd1 vccd1 vccd1 _19194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11043__B1 _09223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18145_ _19835_/Q _18148_/C _18126_/X vssd1 vssd1 vccd1 vccd1 _18145_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_102_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15357_ _15357_/A vssd1 vssd1 vccd1 vccd1 _18727_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14780__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12569_ _12658_/A _12715_/B _15242_/C _12568_/X vssd1 vssd1 vccd1 vccd1 _13440_/S
+ sky130_fd_sc_hd__or4b_2
XANTENNA__14780__B2 _14732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09882__S1 _09881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14308_ _14310_/B _14308_/B vssd1 vssd1 vccd1 vccd1 _14312_/B sky130_fd_sc_hd__and2_1
XANTENNA__09448__S _09448_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18076_ _18075_/A _18075_/C _19812_/Q vssd1 vssd1 vccd1 vccd1 _18077_/C sky130_fd_sc_hd__a21oi_1
XFILLER_8_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15288_ _15288_/A vssd1 vssd1 vccd1 vccd1 _18697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17027_ _17049_/A vssd1 vssd1 vccd1 vccd1 _17036_/S sky130_fd_sc_hd__buf_2
XFILLER_144_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15974__A _16031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14239_ _14059_/A _14241_/B _13975_/A _14238_/X vssd1 vssd1 vccd1 vccd1 _14239_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12543__B1 _12742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15185__S _15185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09780_ _10094_/A vssd1 vssd1 vccd1 vccd1 _10114_/S sky130_fd_sc_hd__buf_2
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18978_ _18982_/CLK _18978_/D vssd1 vssd1 vccd1 vccd1 _18978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _17948_/A _17934_/C vssd1 vssd1 vccd1 vccd1 _17929_/Y sky130_fd_sc_hd__nor2_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15913__S _15913_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09212__A _09212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09214_ _09214_/A vssd1 vssd1 vccd1 vccd1 _09215_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09145_ _09145_/A vssd1 vssd1 vccd1 vccd1 _09146_/A sky130_fd_sc_hd__buf_2
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17575__S _17579_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11189__A _11189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10093__A _10093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_opt_1_0_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__A1 _09927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09950__B2 _18449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09978_ _09978_/A vssd1 vssd1 vccd1 vccd1 _09979_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10821__A _19694_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_133_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12837__A1 _12840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17225__A0 _18451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09702__A1 _09172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11940_ _11940_/A _12030_/A vssd1 vssd1 vccd1 vccd1 _11947_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _11871_/A _11871_/B vssd1 vssd1 vccd1 vccd1 _11872_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10967__S _11027_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12748__A _12748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _13765_/S vssd1 vssd1 vccd1 vccd1 _13758_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_55_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ _10830_/A _10818_/X _10820_/X _10821_/X vssd1 vssd1 vccd1 vccd1 _10823_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _18553_/Q _14577_/X _14589_/X _14585_/X vssd1 vssd1 vccd1 vccd1 _18553_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13541_ _14577_/A _11552_/A _13537_/X _18419_/Q vssd1 vssd1 vccd1 vccd1 _13542_/B
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_1_1_1_clock clkbuf_1_1_1_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_10753_ _18823_/Q _19377_/Q _19539_/Q _18791_/Q _10858_/A _10740_/X vssd1 vssd1 vccd1
+ vccd1 _10753_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14963__A _16709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16260_ _16099_/X _19103_/Q _16268_/S vssd1 vssd1 vccd1 vccd1 _16261_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ _13472_/A vssd1 vssd1 vccd1 vccd1 _18395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10684_ _19636_/Q _19053_/Q _19090_/Q _18696_/Q _10860_/S _09139_/A vssd1 vssd1 vccd1
+ vccd1 _10684_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15211_ _18673_/Q _15210_/X _15217_/S vssd1 vssd1 vccd1 vccd1 _15212_/A sky130_fd_sc_hd__mux2_1
X_12423_ _11202_/A _18520_/Q _12423_/S vssd1 vssd1 vccd1 vccd1 _12424_/A sky130_fd_sc_hd__mux2_8
X_16191_ _16191_/A vssd1 vssd1 vccd1 vccd1 _19068_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12483__A _12483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11120__S0 _10230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15142_ _15142_/A vssd1 vssd1 vccd1 vccd1 _18651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13298__B _18634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12354_ _12354_/A _12354_/B vssd1 vssd1 vccd1 vccd1 _12371_/C sky130_fd_sc_hd__nor2_2
XFILLER_138_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17485__S _17485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11099__A _11099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305_ _11305_/A _14900_/B vssd1 vssd1 vccd1 vccd1 _11381_/C sky130_fd_sc_hd__nand2_2
X_15073_ input25/X _14924_/X _14925_/X vssd1 vssd1 vccd1 vccd1 _15073_/X sky130_fd_sc_hd__a21o_1
XFILLER_142_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12285_ _12285_/A _12285_/B vssd1 vssd1 vccd1 vccd1 _12371_/A sky130_fd_sc_hd__nor2_4
XANTENNA__18170__A _18170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18901_ _19326_/CLK _18901_/D vssd1 vssd1 vccd1 vccd1 _18901_/Q sky130_fd_sc_hd__dfxtp_1
X_14024_ _14026_/A _14026_/B vssd1 vssd1 vccd1 vccd1 _14024_/Y sky130_fd_sc_hd__nand2_1
X_11236_ _11234_/Y _11137_/X _10300_/A _11238_/A vssd1 vssd1 vccd1 vccd1 _11266_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_134_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18832_ _19549_/CLK _18832_/D vssd1 vssd1 vccd1 vccd1 _18832_/Q sky130_fd_sc_hd__dfxtp_1
X_11167_ _19529_/Q _19143_/Q _19593_/Q _18749_/Q _11153_/X _10306_/X vssd1 vssd1 vccd1
+ vccd1 _11168_/B sky130_fd_sc_hd__mux4_1
XFILLER_171_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14203__A _14203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10118_ _10120_/A _10113_/X _10115_/X _10117_/X vssd1 vssd1 vccd1 vccd1 _10118_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_49_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18763_ _19706_/CLK _18763_/D vssd1 vssd1 vccd1 vccd1 _18763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15018__B _15018_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15975_ _14772_/X _18987_/Q _15983_/S vssd1 vssd1 vccd1 vccd1 _15976_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11098_ _19642_/Q _19059_/Q _19096_/Q _18702_/Q _09447_/A _09539_/A vssd1 vssd1 vccd1
+ vccd1 _11099_/B sky130_fd_sc_hd__mux4_1
X_17714_ _17713_/X _12634_/B _17708_/A vssd1 vssd1 vccd1 vccd1 _17714_/X sky130_fd_sc_hd__a21bo_1
XFILLER_36_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10049_ _09892_/X _10042_/X _10044_/X _10048_/X _09395_/X vssd1 vssd1 vccd1 vccd1
+ _10049_/X sky130_fd_sc_hd__a311o_2
X_14926_ input10/X _14924_/X _14925_/X vssd1 vssd1 vccd1 vccd1 _14926_/X sky130_fd_sc_hd__a21o_1
X_18694_ _19636_/CLK _18694_/D vssd1 vssd1 vccd1 vccd1 _18694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17645_ _17645_/A _17649_/C vssd1 vssd1 vccd1 vccd1 _17645_/Y sky130_fd_sc_hd__xnor2_2
X_14857_ _14856_/X _18598_/Q _14880_/S vssd1 vssd1 vccd1 vccd1 _14858_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13808_ _13839_/S _13800_/B _13795_/X _13805_/X _13807_/X vssd1 vssd1 vccd1 vccd1
+ _13808_/X sky130_fd_sc_hd__o221a_1
X_14788_ _18433_/Q _13086_/B _14992_/S vssd1 vssd1 vccd1 vccd1 _14788_/X sky130_fd_sc_hd__mux2_1
X_17576_ _17576_/A vssd1 vssd1 vccd1 vccd1 _19646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19315_ _19541_/CLK _19315_/D vssd1 vssd1 vccd1 vccd1 _19315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16527_ _16573_/S vssd1 vssd1 vccd1 vccd1 _16536_/S sky130_fd_sc_hd__buf_2
X_13739_ _13845_/S vssd1 vssd1 vccd1 vccd1 _13997_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19246_ _19568_/CLK _19246_/D vssd1 vssd1 vccd1 vccd1 _19246_/Q sky130_fd_sc_hd__dfxtp_1
X_16458_ _16071_/X _19190_/Q _16464_/S vssd1 vssd1 vccd1 vccd1 _16459_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15409_ _15409_/A vssd1 vssd1 vccd1 vccd1 _18751_/D sky130_fd_sc_hd__clkbuf_1
X_16389_ _19160_/Q _15532_/X _16391_/S vssd1 vssd1 vccd1 vccd1 _16390_/A sky130_fd_sc_hd__mux2_1
X_19177_ _19595_/CLK _19177_/D vssd1 vssd1 vccd1 vccd1 _19177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10906__A _10906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18128_ _18131_/B _18131_/C _18127_/Y vssd1 vssd1 vccd1 vccd1 _19829_/D sky130_fd_sc_hd__o21a_1
XFILLER_117_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10775__C1 _10774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18059_ _18059_/A _19806_/Q _18059_/C vssd1 vssd1 vccd1 vccd1 _18061_/B sky130_fd_sc_hd__and3_1
X_09901_ _09901_/A _09901_/B vssd1 vssd1 vccd1 vccd1 _09901_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10527__C1 _09392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12840__B _12840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09832_ _10068_/A vssd1 vssd1 vccd1 vccd1 _10044_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09763_ _09763_/A vssd1 vssd1 vccd1 vccd1 _09763_/X sky130_fd_sc_hd__buf_2
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15643__S _15647_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09694_ _11168_/A _09694_/B vssd1 vssd1 vccd1 vccd1 _09694_/X sky130_fd_sc_hd__or2_1
XFILLER_55_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09641__S _10417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09791__S0 _09760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12568__A _14562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14992__A1 _12778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17930__A1 _19761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12755__B1 _12745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09128_ _11376_/A _11484_/A _11374_/A _11296_/C vssd1 vssd1 vccd1 vccd1 _13568_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17694__A0 _12559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16503__A _16503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12070_ _12066_/Y _12069_/X _12165_/S vssd1 vssd1 vccd1 vccd1 _12070_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10518__C1 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16249__A1 _19098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11021_ _09407_/A _11014_/X _11016_/X _11020_/X _09390_/A vssd1 vssd1 vccd1 vccd1
+ _11021_/X sky130_fd_sc_hd__a311o_1
XANTENNA__09923__B2 _18449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11730__A1 _15262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14958__A _14958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15760_ _15806_/S vssd1 vssd1 vccd1 vccd1 _15769_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_46_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _12972_/A _12972_/B _18305_/Q vssd1 vssd1 vccd1 vccd1 _12973_/C sky130_fd_sc_hd__and3_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input11_A io_dbus_rdata[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10297__A1 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11923_ _11871_/A _11921_/Y _11922_/Y vssd1 vssd1 vccd1 vccd1 _11923_/Y sky130_fd_sc_hd__a21oi_1
X_14711_ _14842_/A vssd1 vssd1 vccd1 vccd1 _14711_/X sky130_fd_sc_hd__buf_4
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15691_ _18860_/Q _15526_/X _15697_/S vssd1 vssd1 vccd1 vccd1 _15692_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17430_ _17430_/A vssd1 vssd1 vccd1 vccd1 _19581_/D sky130_fd_sc_hd__clkbuf_1
X_14642_ _14672_/A _14642_/B vssd1 vssd1 vccd1 vccd1 _18567_/D sky130_fd_sc_hd__nor2_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ _11847_/X _11852_/X _11853_/X _12696_/A vssd1 vssd1 vccd1 vccd1 _11854_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12038__A2 _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10049__A1 _09892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10805_ _10805_/A vssd1 vssd1 vccd1 vccd1 _10932_/S sky130_fd_sc_hd__buf_4
X_14573_ _14585_/A vssd1 vssd1 vccd1 vccd1 _14573_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14983__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17361_ _16803_/X _19551_/Q _17363_/S vssd1 vssd1 vccd1 vccd1 _17362_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11785_ _11785_/A _13925_/B vssd1 vssd1 vccd1 vccd1 _11785_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19100_ _19614_/CLK _19100_/D vssd1 vssd1 vccd1 vccd1 _19100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16312_ _16071_/X _19126_/Q _16318_/S vssd1 vssd1 vccd1 vccd1 _16313_/A sky130_fd_sc_hd__mux2_1
X_13524_ _14566_/A _13524_/B _13524_/C _13524_/D vssd1 vssd1 vccd1 vccd1 _13524_/X
+ sky130_fd_sc_hd__or4_1
X_17292_ _17292_/A vssd1 vssd1 vccd1 vccd1 _19520_/D sky130_fd_sc_hd__clkbuf_1
X_10736_ _19313_/Q vssd1 vssd1 vccd1 vccd1 _10736_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16243_ _16243_/A vssd1 vssd1 vccd1 vccd1 _19095_/D sky130_fd_sc_hd__clkbuf_1
X_19031_ _19614_/CLK _19031_/D vssd1 vssd1 vccd1 vccd1 _19031_/Q sky130_fd_sc_hd__dfxtp_1
X_13455_ _13512_/S vssd1 vssd1 vccd1 vccd1 _13464_/S sky130_fd_sc_hd__buf_2
XANTENNA__14735__A1 _18428_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10667_ _10905_/S vssd1 vssd1 vccd1 vccd1 _10668_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__13102__A _17781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12406_ _12406_/A _12406_/B vssd1 vssd1 vccd1 vccd1 _12408_/B sky130_fd_sc_hd__xnor2_4
XFILLER_126_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16174_ _16196_/A vssd1 vssd1 vccd1 vccd1 _16183_/S sky130_fd_sc_hd__buf_2
XFILLER_154_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13386_ _18646_/Q _13386_/B vssd1 vssd1 vccd1 vccd1 _13386_/X sky130_fd_sc_hd__or2_1
X_10598_ _09529_/X _10591_/X _10593_/X _10597_/X _09392_/A vssd1 vssd1 vccd1 vccd1
+ _10598_/X sky130_fd_sc_hd__a311o_1
XANTENNA__15728__S _15730_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15125_ _15125_/A vssd1 vssd1 vccd1 vccd1 _15125_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12337_ _12333_/X _12336_/Y _12452_/S vssd1 vssd1 vccd1 vccd1 _12337_/X sky130_fd_sc_hd__mux2_1
Xoutput108 _13578_/A vssd1 vssd1 vccd1 vccd1 io_dbus_rd_en sky130_fd_sc_hd__buf_2
XFILLER_154_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17509__A _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput119 _12486_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[17] sky130_fd_sc_hd__buf_2
XFILLER_141_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09726__S _10125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15056_ _15055_/X _18615_/Q _15056_/S vssd1 vssd1 vccd1 vccd1 _15057_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15160__A1 _15159_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12268_ _12268_/A _12292_/B vssd1 vssd1 vccd1 vccd1 _12268_/Y sky130_fd_sc_hd__nor2_1
X_14007_ _14005_/B _13658_/X _13714_/X vssd1 vssd1 vccd1 vccd1 _14007_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_96_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11219_ _11205_/Y _11284_/B _11203_/A _11204_/Y vssd1 vssd1 vccd1 vccd1 _11219_/X
+ sky130_fd_sc_hd__a211o_1
X_19864_ _19872_/CLK _19864_/D vssd1 vssd1 vccd1 vccd1 _19864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10461__A _10461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ _13322_/A _12222_/C vssd1 vssd1 vccd1 vccd1 _12199_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput90 _12313_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[25] sky130_fd_sc_hd__buf_2
X_18815_ _19709_/CLK _18815_/D vssd1 vssd1 vccd1 vccd1 _18815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19795_ _19795_/CLK _19795_/D vssd1 vssd1 vccd1 vccd1 _19795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18746_ _19556_/CLK _18746_/D vssd1 vssd1 vccd1 vccd1 _18746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15958_ _17774_/A _15958_/B vssd1 vssd1 vccd1 vccd1 _18980_/D sky130_fd_sc_hd__nor2_2
XFILLER_76_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14909_ _14908_/X _18602_/Q _14941_/S vssd1 vssd1 vccd1 vccd1 _14910_/A sky130_fd_sc_hd__mux2_1
X_18677_ _19590_/CLK _18677_/D vssd1 vssd1 vccd1 vccd1 _18677_/Q sky130_fd_sc_hd__dfxtp_1
X_15889_ _14753_/X _18948_/Q _15891_/S vssd1 vssd1 vccd1 vccd1 _15890_/A sky130_fd_sc_hd__mux2_1
X_17628_ _13197_/X _17627_/Y _17628_/S vssd1 vssd1 vccd1 vccd1 _17628_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16294__S _16296_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17559_ _17605_/S vssd1 vssd1 vccd1 vccd1 _17568_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__10135__S1 _10331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09697__A _09697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17912__A1 _19759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19229_ _19715_/CLK _19229_/D vssd1 vssd1 vccd1 vccd1 _19229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10636__A _10764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17676__A0 _13279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17853__S _17853_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11173__C1 _09248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09815_ _19621_/Q _19459_/Q _18905_/Q _18675_/Q _09803_/X _09810_/X vssd1 vssd1 vccd1
+ vccd1 _09815_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input3_A io_dbus_rdata[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15373__S _15373_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09746_ _18843_/Q _19397_/Q _19559_/Q _18811_/Q _09734_/X _09595_/A vssd1 vssd1 vccd1
+ vccd1 _09747_/B sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_171_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19571_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_86_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09764__S0 _09760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _10329_/A _09674_/Y _09676_/Y _10288_/A vssd1 vssd1 vccd1 vccd1 _09677_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16993__A _17049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10374__S1 _10349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09516__S0 _10450_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_186_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19285_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10126__S1 _09595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11570_ _11560_/X _11563_/X _12219_/S _11625_/A vssd1 vssd1 vccd1 vccd1 _17855_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10521_ _19639_/Q _19056_/Q _19093_/Q _18699_/Q _10500_/X _10501_/X vssd1 vssd1 vccd1
+ vccd1 _10521_/X sky130_fd_sc_hd__mux4_2
XANTENNA__09400__A _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10546__A _10739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13240_ _13240_/A _13240_/B vssd1 vssd1 vccd1 vccd1 _14813_/B sky130_fd_sc_hd__or2_1
XFILLER_136_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10452_ _10239_/X _10449_/Y _10451_/Y _10496_/A vssd1 vssd1 vccd1 vccd1 _10452_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10203__A1 _10103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13171_ _13171_/A _18623_/Q vssd1 vssd1 vccd1 vccd1 _13171_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10383_ _09276_/A _10373_/X _10382_/X _09283_/A _18440_/Q vssd1 vssd1 vccd1 vccd1
+ _10412_/A sky130_fd_sc_hd__a32o_4
XFILLER_151_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12122_ _13312_/A _12123_/C _18367_/Q vssd1 vssd1 vccd1 vccd1 _12122_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09546__S _09793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input59_A io_ibus_inst[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_124_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19680_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12053_ _12067_/B _11928_/X _12048_/Y _12052_/X vssd1 vssd1 vccd1 vccd1 _17882_/B
+ sky130_fd_sc_hd__o22a_1
X_16930_ _16930_/A vssd1 vssd1 vccd1 vccd1 _19374_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11164__C1 _09134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10506__A2 _10494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12900__B1 _12869_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ _18587_/Q _19276_/Q _11051_/S vssd1 vssd1 vccd1 vccd1 _11004_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16861_ _19344_/Q _16657_/X _16869_/S vssd1 vssd1 vccd1 vccd1 _16862_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18600_ _19513_/CLK _18600_/D vssd1 vssd1 vccd1 vccd1 _18600_/Q sky130_fd_sc_hd__dfxtp_1
X_15812_ _15812_/A vssd1 vssd1 vccd1 vccd1 _18913_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_139_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19468_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17064__A _17463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19580_ _19580_/CLK _19580_/D vssd1 vssd1 vccd1 vccd1 _19580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13456__A1 _13197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16792_ _16792_/A vssd1 vssd1 vccd1 vccd1 _19321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18531_ _18618_/CLK _18531_/D vssd1 vssd1 vccd1 vccd1 _18531_/Q sky130_fd_sc_hd__dfxtp_1
X_12955_ _18295_/Q _12957_/C _12954_/Y vssd1 vssd1 vccd1 vccd1 _18295_/D sky130_fd_sc_hd__a21oi_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15743_ _14740_/X _18883_/Q _15747_/S vssd1 vssd1 vccd1 vccd1 _15744_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14200__B _14203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ _18359_/Q vssd1 vssd1 vccd1 vccd1 _13246_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18462_ _18623_/CLK _18462_/D vssd1 vssd1 vccd1 vccd1 _18462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12886_ _12895_/D vssd1 vssd1 vccd1 vccd1 _12893_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _15674_/A vssd1 vssd1 vccd1 vccd1 _18852_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _16774_/X _19574_/Q _17413_/S vssd1 vssd1 vccd1 vccd1 _17414_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11219__B1 _11203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14625_ _14625_/A vssd1 vssd1 vccd1 vccd1 _18562_/D sky130_fd_sc_hd__clkbuf_1
X_11837_ _13653_/A _13984_/A _11837_/C _13996_/A vssd1 vssd1 vccd1 vccd1 _11939_/B
+ sky130_fd_sc_hd__or4b_2
X_18393_ _19687_/CLK _18393_/D vssd1 vssd1 vccd1 vccd1 _18393_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17003__S _17003_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _18539_/Q _14550_/X _14555_/X _14548_/X vssd1 vssd1 vccd1 vccd1 _18539_/D
+ sky130_fd_sc_hd__o211a_1
X_17344_ _16777_/X _19543_/Q _17352_/S vssd1 vssd1 vccd1 vccd1 _17345_/A sky130_fd_sc_hd__mux2_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _11768_/A _11768_/B vssd1 vssd1 vccd1 vccd1 _11768_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13507_ _13507_/A vssd1 vssd1 vccd1 vccd1 _18411_/D sky130_fd_sc_hd__clkbuf_1
X_10719_ _10724_/A vssd1 vssd1 vccd1 vccd1 _10719_/X sky130_fd_sc_hd__buf_6
XFILLER_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17275_ _17275_/A vssd1 vssd1 vccd1 vccd1 _19512_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16842__S _16845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14487_ _18514_/Q _19752_/Q _14487_/S vssd1 vssd1 vccd1 vccd1 _14488_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11699_ _11699_/A _13667_/A vssd1 vssd1 vccd1 vccd1 _11700_/B sky130_fd_sc_hd__nor2_1
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19014_ _19632_/CLK _19014_/D vssd1 vssd1 vccd1 vccd1 _19014_/Q sky130_fd_sc_hd__dfxtp_1
X_13438_ _18381_/Q _13438_/B vssd1 vssd1 vccd1 vccd1 _13438_/X sky130_fd_sc_hd__or2_1
XFILLER_146_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16226_ _16283_/S vssd1 vssd1 vccd1 vccd1 _16235_/S sky130_fd_sc_hd__buf_2
XANTENNA__17658__A0 _13259_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16157_ _16058_/X _19053_/Q _16161_/S vssd1 vssd1 vccd1 vccd1 _16158_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13369_ _18293_/Q _12638_/X _13119_/C _18376_/Q vssd1 vssd1 vccd1 vccd1 _13369_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12671__A _12671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11942__A1 _11511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15108_ _18632_/Q _15102_/X _15104_/X _11130_/A vssd1 vssd1 vccd1 vccd1 _18632_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16088_ _16087_/X _19030_/Q _16097_/S vssd1 vssd1 vccd1 vccd1 _16089_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15039_ _15049_/B _15038_/Y _14737_/A vssd1 vssd1 vccd1 vccd1 _15039_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_142_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19847_ _19851_/CLK _19847_/D vssd1 vssd1 vccd1 vccd1 _19847_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_110_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09600_ _09600_/A vssd1 vssd1 vccd1 vccd1 _09734_/A sky130_fd_sc_hd__buf_2
XFILLER_95_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19778_ _19779_/CLK _19778_/D vssd1 vssd1 vccd1 vccd1 _19778_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13447__A1 _13149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09531_ _09411_/A _09521_/Y _09524_/Y _09527_/Y _09530_/Y vssd1 vssd1 vccd1 vccd1
+ _09531_/X sky130_fd_sc_hd__o32a_1
XANTENNA__09746__S0 _09734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18729_ _19571_/CLK _18729_/D vssd1 vssd1 vccd1 vccd1 _18729_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10356__S1 _09142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09462_ _19659_/Q _19076_/Q _19113_/Q _18719_/Q _10350_/S _09442_/X vssd1 vssd1 vccd1
+ vccd1 _09463_/B sky130_fd_sc_hd__mux4_1
XFILLER_25_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14947__A1 _18446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09393_ _09393_/A vssd1 vssd1 vccd1 vccd1 _09394_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10108__S1 _10103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12565__B _13108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10366__A _10366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_41_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19271_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17149__A _17762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12581__A _12603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15124__B2 _11148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13686__A1 _14138_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_56_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19003_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_87_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11697__A0 _11696_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16199__S _16205_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10595__S1 _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17821__A0 _15191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09737__S0 _09734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09729_ _18612_/Q _19301_/Q _09729_/S vssd1 vssd1 vccd1 vccd1 _09730_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09657__A3 _09656_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12740_ _18299_/Q _13108_/A _13115_/A _18373_/Q _12739_/X vssd1 vssd1 vccd1 vccd1
+ _12740_/X sky130_fd_sc_hd__a221o_1
XFILLER_15_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12671_ _12671_/A vssd1 vssd1 vccd1 vccd1 _12671_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12949__B1 _12948_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14990_/A _18514_/Q _14410_/S vssd1 vssd1 vccd1 vccd1 _14411_/A sky130_fd_sc_hd__mux2_1
X_11622_ _11622_/A _11622_/B _13671_/A vssd1 vssd1 vccd1 vccd1 _11623_/B sky130_fd_sc_hd__or3_1
XFILLER_63_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15390_ _15390_/A vssd1 vssd1 vccd1 vccd1 _18742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09130__A _10823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14341_ _18458_/Q _18490_/Q _14352_/S vssd1 vssd1 vccd1 vccd1 _14342_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11621__B1 _13671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11553_ _15018_/A _11552_/X _14032_/S vssd1 vssd1 vccd1 vccd1 _11554_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16662__S _16671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09290__A1 _15339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10504_ _10498_/A _10499_/X _10503_/X _09681_/A vssd1 vssd1 vccd1 vccd1 _10504_/X
+ sky130_fd_sc_hd__o211a_1
X_17060_ _19433_/Q _16737_/X _17062_/S vssd1 vssd1 vccd1 vccd1 _17061_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14166__A2 _14168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14272_ _14274_/B _14272_/B vssd1 vssd1 vccd1 vccd1 _14276_/B sky130_fd_sc_hd__and2_1
XFILLER_144_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11484_ _11484_/A _11484_/B vssd1 vssd1 vccd1 vccd1 _11485_/A sky130_fd_sc_hd__nand2_2
X_16011_ _16011_/A vssd1 vssd1 vccd1 vccd1 _19003_/D sky130_fd_sc_hd__clkbuf_1
X_13223_ _18275_/Q _13156_/A _12641_/A _13222_/X vssd1 vssd1 vccd1 vccd1 _13223_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__13374__B1 _13369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15278__S _15278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10435_ _10428_/X _10430_/X _10432_/X _10434_/X _09246_/A vssd1 vssd1 vccd1 vccd1
+ _10435_/X sky130_fd_sc_hd__a221o_4
XFILLER_171_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_7_0_clock clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
X_13154_ _18385_/Q _13154_/B vssd1 vssd1 vccd1 vccd1 _13154_/X sky130_fd_sc_hd__and2_1
XANTENNA__10283__S0 _10224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10366_ _10366_/A vssd1 vssd1 vccd1 vccd1 _10367_/A sky130_fd_sc_hd__buf_2
XANTENNA__15115__B2 _10196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output165_A _17909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _12105_/A _12105_/B vssd1 vssd1 vccd1 vccd1 _14168_/A sky130_fd_sc_hd__nand2_4
XFILLER_112_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _19771_/Q _17963_/C _19772_/Q vssd1 vssd1 vccd1 vccd1 _17964_/B sky130_fd_sc_hd__a21oi_1
X_13085_ _18043_/A _12518_/A _12602_/A _12993_/A _13084_/X vssd1 vssd1 vccd1 vccd1
+ _13086_/B sky130_fd_sc_hd__a221o_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10297_ _09428_/A _10286_/X _10295_/X _09625_/A _10296_/Y vssd1 vssd1 vccd1 vccd1
+ _12485_/A sky130_fd_sc_hd__o32a_4
XANTENNA__14874__B1 _14873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19701_ _19703_/CLK _19701_/D vssd1 vssd1 vccd1 vccd1 _19701_/Q sky130_fd_sc_hd__dfxtp_1
X_12036_ _12036_/A _12036_/B vssd1 vssd1 vccd1 vccd1 _12040_/A sky130_fd_sc_hd__nor2_2
X_16913_ _19368_/Q _16734_/X _16913_/S vssd1 vssd1 vccd1 vccd1 _16914_/A sky130_fd_sc_hd__mux2_1
X_17893_ _17909_/A _17893_/B vssd1 vssd1 vccd1 vccd1 _17894_/A sky130_fd_sc_hd__and2_1
XFILLER_66_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10586__S1 _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09750__C1 _09403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19632_ _19632_/CLK _19632_/D vssd1 vssd1 vccd1 vccd1 _19632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16844_ _16844_/A vssd1 vssd1 vccd1 vccd1 _16844_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_181_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14211__A _14211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19563_ _19709_/CLK _19563_/D vssd1 vssd1 vccd1 vccd1 _19563_/Q sky130_fd_sc_hd__dfxtp_1
X_16775_ _16774_/X _19316_/Q _16775_/S vssd1 vssd1 vccd1 vccd1 _16776_/A sky130_fd_sc_hd__mux2_1
X_13987_ _13971_/X _13973_/Y _13986_/X vssd1 vssd1 vccd1 vccd1 _13987_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15741__S _15747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18514_ _18519_/CLK _18514_/D vssd1 vssd1 vccd1 vccd1 _18514_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15726_ _18876_/Q _15577_/X _15730_/S vssd1 vssd1 vccd1 vccd1 _15727_/A sky130_fd_sc_hd__mux2_1
X_12938_ _18289_/Q _12939_/C _18290_/Q vssd1 vssd1 vccd1 vccd1 _12940_/B sky130_fd_sc_hd__a21oi_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19494_ _19786_/CLK _19494_/D vssd1 vssd1 vccd1 vccd1 _19494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18445_ _19695_/CLK _18445_/D vssd1 vssd1 vccd1 vccd1 _18445_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15657_ _15657_/A vssd1 vssd1 vccd1 vccd1 _18845_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15051__A0 _18455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12869_ _18173_/A vssd1 vssd1 vccd1 vccd1 _12869_/X sky130_fd_sc_hd__buf_2
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14608_ _14624_/A _14608_/B vssd1 vssd1 vccd1 vccd1 _14609_/A sky130_fd_sc_hd__and2_1
XFILLER_159_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18376_ _19690_/CLK _18376_/D vssd1 vssd1 vccd1 vccd1 _18376_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_105_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15588_ _15588_/A vssd1 vssd1 vccd1 vccd1 _18815_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11612__A0 _18575_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17327_ _17327_/A vssd1 vssd1 vccd1 vccd1 _19535_/D sky130_fd_sc_hd__clkbuf_1
X_14539_ _18564_/Q _12763_/X _14538_/Y _14535_/X vssd1 vssd1 vccd1 vccd1 _18532_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10186__A _10186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15354__A1 _15155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17258_ _19505_/Q _16654_/X _17258_/S vssd1 vssd1 vccd1 vccd1 _17259_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16209_ _16134_/X _19077_/Q _16209_/S vssd1 vssd1 vccd1 vccd1 _16210_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17189_ _19483_/Q _17188_/X _17189_/S vssd1 vssd1 vccd1 vccd1 _17190_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10179__B1 _09616_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15106__A1 _18630_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15106__B2 _11082_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15916__S _15924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17803__A0 _15165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09741__C1 _09395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10351__B1 _10475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09514_ _09514_/A vssd1 vssd1 vccd1 vccd1 _09515_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18247__B _18247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09445_ _09629_/A vssd1 vssd1 vccd1 vccd1 _09449_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10654__A1 _19187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12576__A _12600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09376_ _10950_/A vssd1 vssd1 vccd1 vccd1 _10762_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16482__S _16486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14791__A _16664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10220_ _10227_/A vssd1 vssd1 vccd1 vccd1 _10447_/A sky130_fd_sc_hd__buf_2
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10151_ _19261_/Q _19032_/Q _18963_/Q _19357_/Q _10154_/S _09146_/A vssd1 vssd1 vccd1
+ vccd1 _10152_/B sky130_fd_sc_hd__mux4_1
XFILLER_106_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14730__S _14762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ _10212_/A _10082_/B vssd1 vssd1 vccd1 vccd1 _10082_/X sky130_fd_sc_hd__or2_1
XFILLER_59_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13910_ _13738_/X _13892_/X _13908_/X _13909_/X vssd1 vssd1 vccd1 vccd1 _13910_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_87_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14890_ _15010_/A vssd1 vssd1 vccd1 vccd1 _14941_/S sky130_fd_sc_hd__buf_4
XFILLER_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13841_ _13839_/X _13840_/X _13881_/S vssd1 vssd1 vccd1 vccd1 _13841_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14084__A1 _18437_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16560_ _16560_/A vssd1 vssd1 vccd1 vccd1 _16569_/S sky130_fd_sc_hd__buf_4
X_13772_ _13637_/X _13631_/X _13775_/S vssd1 vssd1 vccd1 vccd1 _13772_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10984_ _09168_/A _10983_/X _09177_/A vssd1 vssd1 vccd1 vccd1 _10984_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15511_ _18791_/Q _15510_/X _15520_/S vssd1 vssd1 vccd1 vccd1 _15512_/A sky130_fd_sc_hd__mux2_1
X_12723_ _19772_/Q _12629_/S _12722_/X vssd1 vssd1 vccd1 vccd1 _12723_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16491_ _16119_/X _19205_/Q _16497_/S vssd1 vssd1 vccd1 vccd1 _16492_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12486__A _12486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18230_ _18230_/A _18230_/B vssd1 vssd1 vccd1 vccd1 _19864_/D sky130_fd_sc_hd__nor2_1
X_12654_ _18639_/Q _14946_/B _14946_/C _14946_/D vssd1 vssd1 vccd1 vccd1 _12654_/X
+ sky130_fd_sc_hd__or4_1
X_15442_ _18764_/Q _15175_/X _15448_/S vssd1 vssd1 vccd1 vccd1 _15443_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09799__C1 _09231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17488__S _17496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11605_ _14547_/A _11213_/X _11216_/X vssd1 vssd1 vccd1 vccd1 _13585_/B sky130_fd_sc_hd__o21bai_2
X_18161_ _19841_/Q _18164_/C _18126_/X vssd1 vssd1 vccd1 vccd1 _18161_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12585_ _12585_/A vssd1 vssd1 vccd1 vccd1 _12606_/A sky130_fd_sc_hd__buf_2
X_15373_ _18735_/Q _15184_/X _15373_/S vssd1 vssd1 vccd1 vccd1 _15374_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18173__A _18173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_128_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17112_ _17112_/A vssd1 vssd1 vccd1 vccd1 _19455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09795__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14324_ _14324_/A _14324_/B vssd1 vssd1 vccd1 vccd1 _14324_/X sky130_fd_sc_hd__or2_1
XANTENNA__14139__A2 _14138_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11536_ _09113_/B _11474_/B _11339_/X vssd1 vssd1 vccd1 vccd1 _11537_/D sky130_fd_sc_hd__o21a_1
X_18092_ _18094_/A _18094_/C _18082_/X vssd1 vssd1 vccd1 vccd1 _18092_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12933__B _18287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17043_ _19425_/Q _16712_/X _17047_/S vssd1 vssd1 vccd1 vccd1 _17044_/A sky130_fd_sc_hd__mux2_1
X_14255_ _14003_/X _14252_/Y _14254_/X vssd1 vssd1 vccd1 vccd1 _14255_/Y sky130_fd_sc_hd__o21ai_1
X_11467_ _11692_/A vssd1 vssd1 vccd1 vccd1 _11470_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10734__A _10996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13110__A _13110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13206_ _19665_/Q _12668_/X _15242_/D _18389_/Q vssd1 vssd1 vccd1 vccd1 _13206_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10418_ _18861_/Q _19319_/Q _10465_/S vssd1 vssd1 vccd1 vccd1 _10418_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14186_ _18444_/Q _14185_/Y _14209_/S vssd1 vssd1 vccd1 vccd1 _14187_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11398_ _18548_/Q _18547_/Q _18546_/Q _18549_/Q vssd1 vssd1 vccd1 vccd1 _11401_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_98_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13137_ _13183_/B _13136_/X _14673_/A vssd1 vssd1 vccd1 vccd1 _13137_/X sky130_fd_sc_hd__a21o_1
XFILLER_124_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10349_ _10349_/A _10349_/B vssd1 vssd1 vccd1 vccd1 _10349_/X sky130_fd_sc_hd__and2_1
X_18994_ _19223_/CLK _18994_/D vssd1 vssd1 vccd1 vccd1 _18994_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10008__S0 _10075_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17945_ _17980_/A _17945_/B _17945_/C vssd1 vssd1 vccd1 vccd1 _19766_/D sky130_fd_sc_hd__nor3_1
X_13068_ _17935_/A _13068_/B _13068_/C vssd1 vssd1 vccd1 vccd1 _18332_/D sky130_fd_sc_hd__nor3_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12019_ _13265_/A _12020_/C _18363_/Q vssd1 vssd1 vccd1 vccd1 _12019_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17876_ _17882_/A _17876_/B vssd1 vssd1 vccd1 vccd1 _17877_/A sky130_fd_sc_hd__or2_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19615_ _19647_/CLK _19615_/D vssd1 vssd1 vccd1 vccd1 _19615_/Q sky130_fd_sc_hd__dfxtp_1
X_16827_ _16825_/X _19332_/Q _16839_/S vssd1 vssd1 vccd1 vccd1 _16828_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16567__S _16569_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19546_ _19546_/CLK _19546_/D vssd1 vssd1 vccd1 vccd1 _19546_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13283__C1 _13282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16758_ _16758_/A vssd1 vssd1 vccd1 vccd1 _16758_/X sky130_fd_sc_hd__buf_2
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10097__C1 _09249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15709_ _15709_/A vssd1 vssd1 vccd1 vccd1 _18868_/D sky130_fd_sc_hd__clkbuf_1
X_19477_ _19488_/CLK _19477_/D vssd1 vssd1 vccd1 vccd1 _19477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16689_ _16689_/A vssd1 vssd1 vccd1 vccd1 _16689_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09230_ _09230_/A vssd1 vssd1 vccd1 vccd1 _09231_/A sky130_fd_sc_hd__clkbuf_4
X_18428_ _19078_/CLK _18428_/D vssd1 vssd1 vccd1 vccd1 _18428_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16772__A0 _16771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09161_ _10011_/S vssd1 vssd1 vccd1 vccd1 _09911_/S sky130_fd_sc_hd__buf_2
XANTENNA__17398__S _17402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18359_ _19082_/CLK _18359_/D vssd1 vssd1 vccd1 vccd1 _18359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10495__S0 _10242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09092_ _09125_/A _18566_/Q vssd1 vssd1 vccd1 vccd1 _11313_/D sky130_fd_sc_hd__or2_2
XFILLER_147_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12474__A_N _12472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10247__S0 _11110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09994_ _09908_/A _09993_/X _10007_/A vssd1 vssd1 vccd1 vccd1 _09994_/X sky130_fd_sc_hd__o21a_1
XFILLER_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10979__A1_N _12462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11922__B _13614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09428_ _09428_/A vssd1 vssd1 vccd1 vccd1 _09429_/A sky130_fd_sc_hd__buf_2
XANTENNA__16763__A0 _16761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11435__C_N _18417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09359_ _11189_/A vssd1 vssd1 vccd1 vccd1 _10132_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12370_ _12361_/A _12186_/X _12365_/X _12369_/X vssd1 vssd1 vccd1 vccd1 _12370_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11321_ _18585_/Q _11321_/B _11321_/C vssd1 vssd1 vccd1 vccd1 _11322_/D sky130_fd_sc_hd__and3b_1
XFILLER_153_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14040_ _14040_/A vssd1 vssd1 vccd1 vccd1 _14040_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11252_ _11252_/A _10881_/X vssd1 vssd1 vccd1 vccd1 _11254_/B sky130_fd_sc_hd__or2b_1
XFILLER_141_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15556__S _15568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ _10103_/X _10200_/X _10202_/X vssd1 vssd1 vccd1 vccd1 _10203_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11183_ _09616_/X _11176_/Y _11178_/Y _11180_/Y _11182_/Y vssd1 vssd1 vccd1 vccd1
+ _11183_/X sky130_fd_sc_hd__o32a_1
XFILLER_121_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input41_A io_ibus_inst[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ _18772_/Q _19001_/Q _18932_/Q _19230_/Q _10125_/X _09595_/A vssd1 vssd1 vccd1
+ vccd1 _10134_/X sky130_fd_sc_hd__mux4_1
X_15991_ _15991_/A vssd1 vssd1 vccd1 vccd1 _18994_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17730_ _17730_/A vssd1 vssd1 vccd1 vccd1 _17730_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10065_ _19649_/Q _19066_/Q _19103_/Q _18709_/Q _09808_/A _09936_/A vssd1 vssd1 vccd1
+ vccd1 _10065_/X sky130_fd_sc_hd__mux4_1
X_14942_ _14942_/A vssd1 vssd1 vccd1 vccd1 _18605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_54_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17661_ _17661_/A vssd1 vssd1 vccd1 vccd1 _19669_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09720__A2 _09710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14873_ _14873_/A _14873_/B _14873_/C _14873_/D vssd1 vssd1 vccd1 vccd1 _14873_/X
+ sky130_fd_sc_hd__or4_2
XANTENNA__16387__S _16391_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19400_ _19624_/CLK _19400_/D vssd1 vssd1 vccd1 vccd1 _19400_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10961__S1 _10960_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16612_ _16612_/A vssd1 vssd1 vccd1 vccd1 _19261_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12068__B1 _19743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13824_ _13821_/A _13808_/X _13821_/Y _13823_/X vssd1 vssd1 vccd1 vccd1 _13824_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17592_ _17592_/A vssd1 vssd1 vccd1 vccd1 _17601_/S sky130_fd_sc_hd__buf_4
XFILLER_90_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19331_ _19331_/CLK _19331_/D vssd1 vssd1 vccd1 vccd1 _19331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16543_ _19228_/Q _15545_/X _16547_/S vssd1 vssd1 vccd1 vccd1 _16544_/A sky130_fd_sc_hd__mux2_1
X_13755_ _13682_/X _13678_/X _13758_/S vssd1 vssd1 vccd1 vccd1 _13755_/X sky130_fd_sc_hd__mux2_1
X_10967_ _18852_/Q _19310_/Q _11027_/S vssd1 vssd1 vccd1 vccd1 _10967_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12706_ _18301_/Q _12564_/A _13418_/S _19480_/Q _12705_/X vssd1 vssd1 vccd1 vccd1
+ _12706_/X sky130_fd_sc_hd__a221o_1
X_19262_ _19648_/CLK _19262_/D vssd1 vssd1 vccd1 vccd1 _19262_/Q sky130_fd_sc_hd__dfxtp_1
X_16474_ _16474_/A vssd1 vssd1 vccd1 vccd1 _19197_/D sky130_fd_sc_hd__clkbuf_1
X_13686_ _14155_/B _14138_/B _13689_/S vssd1 vssd1 vccd1 vccd1 _13686_/X sky130_fd_sc_hd__mux2_1
X_10898_ _18819_/Q _19373_/Q _19535_/Q _18787_/Q _10648_/S _10785_/X vssd1 vssd1 vccd1
+ vccd1 _10899_/B sky130_fd_sc_hd__mux4_1
X_18213_ _19858_/Q _18210_/A _18212_/Y vssd1 vssd1 vccd1 vccd1 _19858_/D sky130_fd_sc_hd__o21a_1
X_15425_ _15425_/A vssd1 vssd1 vccd1 vccd1 _18756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12637_ _13156_/A vssd1 vssd1 vccd1 vccd1 _13270_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_19193_ _19710_/CLK _19193_/D vssd1 vssd1 vccd1 vccd1 _19193_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12944__A _12991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18144_ _19834_/Q _18141_/C _18143_/Y vssd1 vssd1 vccd1 vccd1 _19834_/D sky130_fd_sc_hd__o21a_1
XFILLER_157_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11043__A1 _10996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09729__S _09729_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12568_ _14562_/A _15242_/B vssd1 vssd1 vccd1 vccd1 _12568_/X sky130_fd_sc_hd__and2_2
XFILLER_145_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15356_ _18727_/Q _15159_/X _15362_/S vssd1 vssd1 vccd1 vccd1 _15357_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14307_ _14307_/A vssd1 vssd1 vccd1 vccd1 _18454_/D sky130_fd_sc_hd__clkbuf_1
X_11519_ _11519_/A _11519_/B _11519_/C _11519_/D vssd1 vssd1 vccd1 vccd1 _11665_/C
+ sky130_fd_sc_hd__or4_1
X_18075_ _18075_/A _19812_/Q _18075_/C vssd1 vssd1 vccd1 vccd1 _18077_/B sky130_fd_sc_hd__and3_1
XFILLER_171_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15287_ _18697_/Q _15165_/X _15289_/S vssd1 vssd1 vccd1 vccd1 _15288_/A sky130_fd_sc_hd__mux2_1
X_12499_ _12499_/A _12503_/B vssd1 vssd1 vccd1 vccd1 _12499_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17026_ _17026_/A vssd1 vssd1 vccd1 vccd1 _19417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14238_ _14262_/A _14241_/A vssd1 vssd1 vccd1 vccd1 _14238_/X sky130_fd_sc_hd__and2_1
XFILLER_172_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15466__S _15470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14169_ _13943_/A _14164_/Y _14168_/Y vssd1 vssd1 vccd1 vccd1 _14169_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__17247__A _17391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _18982_/CLK _18977_/D vssd1 vssd1 vccd1 vccd1 _18977_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _17936_/D vssd1 vssd1 vccd1 vccd1 _17934_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17859_ _11684_/A _11684_/B _14638_/A vssd1 vssd1 vccd1 vccd1 _19730_/D sky130_fd_sc_hd__a21o_1
XFILLER_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18078__A _18199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19529_ _19625_/CLK _19529_/D vssd1 vssd1 vccd1 vccd1 _19529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09570__S1 _09642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09213_ _09689_/A vssd1 vssd1 vccd1 vccd1 _09214_/A sky130_fd_sc_hd__buf_2
XFILLER_167_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09144_ _09144_/A vssd1 vssd1 vccd1 vccd1 _09145_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_147_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12782__A1 _12731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12782__B2 _12763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15376__S _15384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09950__A2 _09940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11917__B _13622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09977_ _10010_/S _09954_/Y _09976_/Y _09763_/A vssd1 vssd1 vccd1 vccd1 _09977_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_58_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_opt_5_0_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17225__A1 _13364_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10312__A3 _19354_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6_0_clock clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_6_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_73_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11870_ _11870_/A _13617_/A vssd1 vssd1 vccd1 vccd1 _11871_/B sky130_fd_sc_hd__or2_1
XFILLER_44_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _19694_/Q vssd1 vssd1 vccd1 vccd1 _10821_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09403__A _09403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11652__B _13665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13262__A2 _13259_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10752_ _10752_/A _10752_/B vssd1 vssd1 vccd1 vccd1 _10752_/X sky130_fd_sc_hd__or2_1
X_13540_ _13540_/A vssd1 vssd1 vccd1 vccd1 _18418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13471_ _18395_/Q _12727_/X _13475_/S vssd1 vssd1 vccd1 vccd1 _13472_/A sky130_fd_sc_hd__mux2_1
X_10683_ _10875_/A _10683_/B vssd1 vssd1 vccd1 vccd1 _10683_/X sky130_fd_sc_hd__or2_1
XFILLER_139_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09218__B2 _09856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15210_ _16712_/A vssd1 vssd1 vccd1 vccd1 _15210_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15140__A _15239_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12422_ _14324_/A _12422_/B vssd1 vssd1 vccd1 vccd1 _12426_/A sky130_fd_sc_hd__xor2_1
XFILLER_139_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16190_ _16106_/X _19068_/Q _16194_/S vssd1 vssd1 vccd1 vccd1 _16191_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11120__S1 _10245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15141_ _18651_/Q _15133_/X _15153_/S vssd1 vssd1 vccd1 vccd1 _15142_/A sky130_fd_sc_hd__mux2_1
X_12353_ _12353_/A _12372_/A vssd1 vssd1 vccd1 vccd1 _12354_/B sky130_fd_sc_hd__and2_1
XANTENNA__17161__A0 _18432_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11304_ _18423_/Q _18422_/Q vssd1 vssd1 vccd1 vccd1 _14900_/B sky130_fd_sc_hd__nor2_2
X_15072_ _15069_/Y _15070_/X _15071_/X _14875_/X vssd1 vssd1 vccd1 vccd1 _15072_/X
+ sky130_fd_sc_hd__o22a_1
X_12284_ _12284_/A _14253_/A vssd1 vssd1 vccd1 vccd1 _12285_/B sky130_fd_sc_hd__nor2_1
X_18900_ _19584_/CLK _18900_/D vssd1 vssd1 vccd1 vccd1 _18900_/Q sky130_fd_sc_hd__dfxtp_1
X_14023_ _14126_/A _14026_/B _14022_/X vssd1 vssd1 vccd1 vccd1 _14023_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13595__A _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11235_ _11235_/A _11239_/A _11235_/C vssd1 vssd1 vccd1 vccd1 _11238_/A sky130_fd_sc_hd__and3_1
XFILLER_4_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18831_ _19223_/CLK _18831_/D vssd1 vssd1 vccd1 vccd1 _18831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11166_ _11166_/A _11166_/B vssd1 vssd1 vccd1 vccd1 _11166_/X sky130_fd_sc_hd__or2_1
XFILLER_150_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10117_ _09979_/X _10116_/X _09996_/A vssd1 vssd1 vccd1 vccd1 _10117_/X sky130_fd_sc_hd__a21o_1
X_18762_ _19541_/CLK _18762_/D vssd1 vssd1 vccd1 vccd1 _18762_/Q sky130_fd_sc_hd__dfxtp_1
X_15974_ _16031_/S vssd1 vssd1 vccd1 vccd1 _15983_/S sky130_fd_sc_hd__buf_2
X_11097_ _11097_/A _11097_/B vssd1 vssd1 vccd1 vccd1 _11097_/X sky130_fd_sc_hd__or2_1
XFILLER_95_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17713_ _17730_/A vssd1 vssd1 vccd1 vccd1 _17713_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10839__A1 _10887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10048_ _09385_/A _10045_/X _10047_/X _09319_/A vssd1 vssd1 vccd1 vccd1 _10048_/X
+ sky130_fd_sc_hd__o211a_1
X_14925_ _14925_/A vssd1 vssd1 vccd1 vccd1 _14925_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18693_ _19700_/CLK _18693_/D vssd1 vssd1 vccd1 vccd1 _18693_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12939__A _18290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11843__A _11843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17006__S _17014_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17644_ _17644_/A vssd1 vssd1 vccd1 vccd1 _19666_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13238__C1 _13237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14856_ _16784_/A vssd1 vssd1 vccd1 vccd1 _14856_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13807_ _13839_/S _13800_/B _13806_/X vssd1 vssd1 vccd1 vccd1 _13807_/X sky130_fd_sc_hd__a21o_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17575_ _19646_/Q _16800_/A _17579_/S vssd1 vssd1 vccd1 vccd1 _17576_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16845__S _16845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14450__A1 _19735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14787_ _14787_/A _14796_/B vssd1 vssd1 vccd1 vccd1 _14787_/Y sky130_fd_sc_hd__nor2_1
X_11999_ _11999_/A vssd1 vssd1 vccd1 vccd1 _12116_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19314_ _19539_/CLK _19314_/D vssd1 vssd1 vccd1 vccd1 _19314_/Q sky130_fd_sc_hd__dfxtp_1
X_16526_ _16526_/A vssd1 vssd1 vccd1 vccd1 _19220_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13738_ _14054_/A vssd1 vssd1 vccd1 vccd1 _13738_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19245_ _19633_/CLK _19245_/D vssd1 vssd1 vccd1 vccd1 _19245_/Q sky130_fd_sc_hd__dfxtp_1
X_16457_ _16457_/A vssd1 vssd1 vccd1 vccd1 _19189_/D sky130_fd_sc_hd__clkbuf_1
X_13669_ _13666_/X _13668_/X _13742_/S vssd1 vssd1 vccd1 vccd1 _13669_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15408_ _18751_/Q _15235_/X _15410_/S vssd1 vssd1 vccd1 vccd1 _15409_/A sky130_fd_sc_hd__mux2_1
X_19176_ _19725_/CLK _19176_/D vssd1 vssd1 vccd1 vccd1 _19176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16388_ _16388_/A vssd1 vssd1 vccd1 vccd1 _19159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12393__B _13388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12764__A1 _12731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18127_ _18131_/B _18131_/C _18126_/X vssd1 vssd1 vccd1 vccd1 _18127_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12764__B2 _12763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15985__A _16031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15339_ _15339_/A _16919_/B _15412_/C vssd1 vssd1 vccd1 vccd1 _17391_/B sky130_fd_sc_hd__or3_4
XFILLER_118_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09983__A _10200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18058_ _18059_/A _18059_/C _18057_/Y vssd1 vssd1 vccd1 vccd1 _19805_/D sky130_fd_sc_hd__o21a_1
XFILLER_105_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10870__S0 _10664_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17009_ _17009_/A vssd1 vssd1 vccd1 vccd1 _19409_/D sky130_fd_sc_hd__clkbuf_1
X_09900_ _09755_/A _09756_/A _11152_/C _09899_/Y vssd1 vssd1 vccd1 vccd1 _09901_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_99_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09831_ _18777_/Q _19006_/Q _18937_/Q _19235_/Q _09928_/A _09875_/A vssd1 vssd1 vccd1
+ vccd1 _09831_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15924__S _15924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _09984_/A vssd1 vssd1 vccd1 vccd1 _09763_/A sky130_fd_sc_hd__buf_2
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09693_ _19269_/Q _19040_/Q _18971_/Q _19365_/Q _10257_/S _09542_/A vssd1 vssd1 vccd1
+ vccd1 _09694_/B sky130_fd_sc_hd__mux4_1
XFILLER_27_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09791__S1 _09763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09223__A _09223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14441__A1 _19731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12452__A0 _12450_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17586__S _17590_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12755__A1 _19847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09127_ _11321_/C _14519_/A _11320_/A vssd1 vssd1 vccd1 vccd1 _11296_/C sky130_fd_sc_hd__and3b_1
XANTENNA__17143__A0 _11022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16503__B _16503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13180__A1 _19828_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ _10807_/A _11017_/X _11019_/X _10728_/A vssd1 vssd1 vccd1 vccd1 _11020_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09923__A2 _09910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11169__S1 _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _12972_/A _12972_/B _18305_/Q vssd1 vssd1 vccd1 vccd1 _12973_/B sky130_fd_sc_hd__a21oi_1
XFILLER_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15135__A _16430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14710_ _14903_/A vssd1 vssd1 vccd1 vccd1 _14842_/A sky130_fd_sc_hd__buf_2
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _11922_/A _13614_/A vssd1 vssd1 vccd1 vccd1 _11922_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10297__A2 _10286_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15690_ _15690_/A vssd1 vssd1 vccd1 vccd1 _18859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12478__B _12478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09133__A _09133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14641_ input38/X _14640_/X _14597_/X _14545_/A vssd1 vssd1 vccd1 vccd1 _14642_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _19666_/Q _11959_/B vssd1 vssd1 vccd1 vccd1 _11853_/X sky130_fd_sc_hd__or2_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14974__A _16712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16665__S _16671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _18821_/Q _19375_/Q _19537_/Q _18789_/Q _10724_/X _10726_/X vssd1 vssd1 vccd1
+ vccd1 _10804_/X sky130_fd_sc_hd__mux4_1
X_17360_ _17360_/A vssd1 vssd1 vccd1 vccd1 _19550_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14572_ _14572_/A _14572_/B vssd1 vssd1 vccd1 vccd1 _14572_/Y sky130_fd_sc_hd__nand2_1
X_11784_ _11784_/A vssd1 vssd1 vccd1 vccd1 _13925_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_82_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16311_ _16311_/A vssd1 vssd1 vccd1 vccd1 _19125_/D sky130_fd_sc_hd__clkbuf_1
X_13523_ _14584_/A _13523_/B _14568_/A _11517_/B vssd1 vssd1 vccd1 vccd1 _13524_/D
+ sky130_fd_sc_hd__or4bb_1
X_17291_ _19520_/Q _16702_/X _17291_/S vssd1 vssd1 vccd1 vccd1 _17292_/A sky130_fd_sc_hd__mux2_1
X_10735_ _10548_/X _10733_/X _10871_/A vssd1 vssd1 vccd1 vccd1 _10735_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_40_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19030_ _19614_/CLK _19030_/D vssd1 vssd1 vccd1 vccd1 _19030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16242_ _16074_/X _19095_/Q _16246_/S vssd1 vssd1 vccd1 vccd1 _16243_/A sky130_fd_sc_hd__mux2_1
X_13454_ _13454_/A vssd1 vssd1 vccd1 vccd1 _18387_/D sky130_fd_sc_hd__clkbuf_1
X_10666_ _19314_/Q vssd1 vssd1 vccd1 vccd1 _10666_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14735__A2 _14958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17496__S _17496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12405_ _12385_/A _12385_/B _12384_/A vssd1 vssd1 vccd1 vccd1 _12406_/B sky130_fd_sc_hd__a21oi_2
X_13385_ hold2/A _13123_/X _13382_/X _13384_/X vssd1 vssd1 vccd1 vccd1 _13386_/B sky130_fd_sc_hd__a211o_1
XFILLER_127_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16173_ _16173_/A vssd1 vssd1 vccd1 vccd1 _19060_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10597_ _10524_/A _10594_/X _10596_/X _09314_/A vssd1 vssd1 vccd1 vccd1 _10597_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_166_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15124_ _18643_/Q _15123_/X _15118_/X _11148_/A vssd1 vssd1 vccd1 vccd1 _18643_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12336_ _12336_/A _12387_/C vssd1 vssd1 vccd1 vccd1 _12336_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10852__S0 _10770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput109 _12495_/B vssd1 vssd1 vccd1 vccd1 io_dbus_st_type[0] sky130_fd_sc_hd__buf_2
XFILLER_115_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11838__A _11940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12267_ _19750_/Q _19751_/Q _12267_/C vssd1 vssd1 vccd1 vccd1 _12292_/B sky130_fd_sc_hd__and3_1
X_15055_ _16838_/A vssd1 vssd1 vccd1 vccd1 _15055_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14214__A _14216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14006_ _13978_/X _13658_/X _13797_/A _14005_/X vssd1 vssd1 vccd1 vccd1 _14006_/X
+ sky130_fd_sc_hd__o211a_1
X_11218_ _13568_/A _11284_/B _11284_/C _11208_/Y _11217_/X vssd1 vssd1 vccd1 vccd1
+ _11565_/A sky130_fd_sc_hd__a311o_1
X_19863_ _19872_/CLK _19863_/D vssd1 vssd1 vccd1 vccd1 _19863_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11557__B _13532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12198_ _13322_/A _12222_/C vssd1 vssd1 vccd1 vccd1 _12198_/X sky130_fd_sc_hd__or2_1
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11182__B1 _09616_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput80 _12096_/B vssd1 vssd1 vccd1 vccd1 io_dbus_addr[16] sky130_fd_sc_hd__buf_2
XANTENNA__10461__B _12480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput91 _12333_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[26] sky130_fd_sc_hd__buf_2
XFILLER_68_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11149_ _11149_/A _11149_/B vssd1 vssd1 vccd1 vccd1 _11225_/A sky130_fd_sc_hd__nor2_1
X_18814_ _19626_/CLK _18814_/D vssd1 vssd1 vccd1 vccd1 _18814_/Q sky130_fd_sc_hd__dfxtp_1
X_19794_ _19795_/CLK _19794_/D vssd1 vssd1 vccd1 vccd1 _19794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18745_ _19427_/CLK _18745_/D vssd1 vssd1 vccd1 vccd1 _18745_/Q sky130_fd_sc_hd__dfxtp_1
X_15957_ _15957_/A vssd1 vssd1 vccd1 vccd1 _18979_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14908_ _16797_/A vssd1 vssd1 vccd1 vccd1 _14908_/X sky130_fd_sc_hd__clkbuf_2
X_18676_ _19622_/CLK _18676_/D vssd1 vssd1 vccd1 vccd1 _18676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15888_ _15888_/A vssd1 vssd1 vccd1 vccd1 _18947_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17627_ _17632_/A _17632_/C vssd1 vssd1 vccd1 vccd1 _17627_/Y sky130_fd_sc_hd__xnor2_4
X_14839_ _18437_/Q _12711_/B _14839_/S vssd1 vssd1 vccd1 vccd1 _14839_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09978__A _09978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17260__A _17317_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17558_ _17558_/A vssd1 vssd1 vccd1 vccd1 _19638_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16509_ _16509_/A vssd1 vssd1 vccd1 vccd1 _19212_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17489_ _17489_/A vssd1 vssd1 vccd1 vccd1 _19607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10917__A _19695_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19228_ _19642_/CLK _19228_/D vssd1 vssd1 vccd1 vccd1 _19228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14108__B _14111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_176_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19159_ _19223_/CLK _19159_/D vssd1 vssd1 vccd1 vccd1 _19159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11096__S0 _10348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10843__S0 _11050_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11748__A _11751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_87_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15654__S _15658_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09814_ _09814_/A _09814_/B vssd1 vssd1 vccd1 vccd1 _09814_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09745_ _10144_/A _09744_/X _09414_/A vssd1 vssd1 vccd1 vccd1 _09745_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_28_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09669__A1 _09412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09764__S1 _09763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09676_ _09735_/A _09676_/B vssd1 vssd1 vccd1 vccd1 _09676_/Y sky130_fd_sc_hd__nand2_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10099__A _12489_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09516__S1 _09587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11930__B _11930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10520_ _10524_/A _10520_/B vssd1 vssd1 vccd1 vccd1 _10520_/X sky130_fd_sc_hd__or2_1
XFILLER_52_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12728__A1 _13106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10451_ _10451_/A _10451_/B vssd1 vssd1 vccd1 vccd1 _10451_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13170_ _18353_/Q _13118_/X _13169_/X vssd1 vssd1 vccd1 vccd1 _18353_/D sky130_fd_sc_hd__a21o_1
X_10382_ _10375_/X _10377_/X _10379_/X _10381_/X _09247_/A vssd1 vssd1 vccd1 vccd1
+ _10382_/X sky130_fd_sc_hd__a221o_4
XFILLER_124_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12121_ _12098_/B _12119_/X _12120_/Y vssd1 vssd1 vccd1 vccd1 _12121_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12052_ _11885_/X _12050_/X _12051_/Y _11625_/A vssd1 vssd1 vccd1 vccd1 _12052_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_151_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11003_ _09480_/A _11003_/B vssd1 vssd1 vccd1 vccd1 _11003_/X sky130_fd_sc_hd__and2b_1
XANTENNA__10506__A3 _10505_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16860_ _16917_/S vssd1 vssd1 vccd1 vccd1 _16869_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15811_ _14714_/X _18913_/Q _15819_/S vssd1 vssd1 vccd1 vccd1 _15812_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13592__B _13724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17064__B _17064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16791_ _16790_/X _19321_/Q _16791_/S vssd1 vssd1 vccd1 vccd1 _16792_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14653__A1 _14555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14653__B2 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18530_ _18618_/CLK _18530_/D vssd1 vssd1 vccd1 vccd1 _18530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15742_ _15742_/A vssd1 vssd1 vccd1 vccd1 _18882_/D sky130_fd_sc_hd__clkbuf_1
X_12954_ _18295_/Q _12957_/C _12948_/X vssd1 vssd1 vccd1 vccd1 _12954_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _11847_/X _11903_/X _11904_/X _12696_/A vssd1 vssd1 vccd1 vccd1 _11905_/X
+ sky130_fd_sc_hd__o211a_1
X_18461_ _18623_/CLK _18461_/D vssd1 vssd1 vccd1 vccd1 _18461_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_clock clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output110_A _13570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15673_ _18852_/Q _15500_/X _15675_/S vssd1 vssd1 vccd1 vccd1 _15674_/A sky130_fd_sc_hd__mux2_1
X_12885_ _18275_/Q _18274_/Q _18273_/Q _12885_/D vssd1 vssd1 vccd1 vccd1 _12895_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__13208__A2 _13130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _17412_/A vssd1 vssd1 vccd1 vccd1 _19573_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _14624_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14625_/A sky130_fd_sc_hd__and2_1
X_18392_ _19496_/CLK _18392_/D vssd1 vssd1 vccd1 vccd1 _18392_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _13761_/A _11836_/B vssd1 vssd1 vccd1 vccd1 _11837_/C sky130_fd_sc_hd__or2_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _17389_/S vssd1 vssd1 vccd1 vccd1 _17352_/S sky130_fd_sc_hd__buf_4
X_14555_ _14555_/A _14559_/B vssd1 vssd1 vccd1 vccd1 _14555_/X sky130_fd_sc_hd__or2_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _11767_/A _11766_/X vssd1 vssd1 vccd1 vccd1 _11768_/B sky130_fd_sc_hd__or2b_1
XANTENNA__10737__A _10982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13506_ _18411_/Q _13399_/X _13508_/S vssd1 vssd1 vccd1 vccd1 _13507_/A sky130_fd_sc_hd__mux2_1
X_17274_ _19512_/Q _16677_/X _17280_/S vssd1 vssd1 vccd1 vccd1 _17275_/A sky130_fd_sc_hd__mux2_1
X_10718_ _10807_/A vssd1 vssd1 vccd1 vccd1 _10946_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14486_ _14486_/A vssd1 vssd1 vccd1 vccd1 _18513_/D sky130_fd_sc_hd__clkbuf_1
X_11698_ _11699_/A _13667_/A vssd1 vssd1 vccd1 vccd1 _11746_/A sky130_fd_sc_hd__and2_1
XANTENNA__12719__A1 _18279_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19013_ _19804_/CLK _19013_/D vssd1 vssd1 vccd1 vccd1 _19013_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15739__S _15747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16225_ _16225_/A vssd1 vssd1 vccd1 vccd1 _19087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13437_ _15262_/B vssd1 vssd1 vccd1 vccd1 _13437_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_146_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12952__A _18294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10649_ _10649_/A vssd1 vssd1 vccd1 vccd1 _10649_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13392__A1 _19687_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17658__A1 _17657_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16156_ _16156_/A vssd1 vssd1 vccd1 vccd1 _19052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13368_ _13403_/A _18645_/Q vssd1 vssd1 vccd1 vccd1 _13368_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11568__A input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15107_ _18631_/Q _15102_/X _15104_/X _10461_/A vssd1 vssd1 vccd1 vccd1 _18631_/D
+ sky130_fd_sc_hd__a22o_1
X_12319_ _13352_/A _12320_/C _18375_/Q vssd1 vssd1 vccd1 vccd1 _12319_/Y sky130_fd_sc_hd__a21oi_1
X_16087_ _16797_/A vssd1 vssd1 vccd1 vccd1 _16087_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13299_ _19871_/Q _12603_/A _12583_/A _19839_/Q vssd1 vssd1 vccd1 vccd1 _13299_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15038_ _15027_/A _15037_/C _18486_/Q vssd1 vssd1 vccd1 vccd1 _15038_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_170_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09443__S0 _10350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14879__A _16790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19846_ _19866_/CLK _19846_/D vssd1 vssd1 vccd1 vccd1 _19846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19777_ _19779_/CLK _19777_/D vssd1 vssd1 vccd1 vccd1 _19777_/Q sky130_fd_sc_hd__dfxtp_1
X_16989_ _16989_/A vssd1 vssd1 vccd1 vccd1 _19401_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12399__A _14310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09530_ _10498_/A _09528_/X _09529_/X vssd1 vssd1 vccd1 vccd1 _09530_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09746__S1 _09595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18728_ _19636_/CLK _18728_/D vssd1 vssd1 vccd1 vccd1 _18728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09461_ _09434_/X _09444_/X _09453_/X _09460_/X _10373_/A vssd1 vssd1 vccd1 vccd1
+ _09461_/X sky130_fd_sc_hd__a311o_2
X_18659_ _19444_/CLK _18659_/D vssd1 vssd1 vccd1 vccd1 _18659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09392_ _09392_/A vssd1 vssd1 vccd1 vccd1 _09393_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10647__A _11050_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17897__A1 _19749_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17149__B _17149_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10816__S0 _10982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15384__S _15384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09985__S1 _09984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09728_ _09728_/A vssd1 vssd1 vccd1 vccd1 _09867_/A sky130_fd_sc_hd__buf_2
XANTENNA__09737__S1 _10186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10657__C1 _09392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ _09671_/A _09659_/B vssd1 vssd1 vccd1 vccd1 _09659_/Y sky130_fd_sc_hd__nor2_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17104__S _17108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11941__A _14589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12541_/C _14562_/A _12670_/C vssd1 vssd1 vccd1 vccd1 _12671_/A sky130_fd_sc_hd__and3b_2
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12756__B _12756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12949__A1 _18293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11622_/A _11622_/B _13671_/A vssd1 vssd1 vccd1 vccd1 _11621_/X sky130_fd_sc_hd__o21a_1
XANTENNA__17337__A0 _16768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14340_ _14384_/A vssd1 vssd1 vccd1 vccd1 _14352_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_129_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11552_ _11552_/A _11552_/B _11551_/Y vssd1 vssd1 vccd1 vccd1 _11552_/X sky130_fd_sc_hd__or3b_2
XFILLER_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15559__S _15568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10503_ _10524_/A _10503_/B vssd1 vssd1 vccd1 vccd1 _10503_/X sky130_fd_sc_hd__or2_1
X_14271_ _18451_/Q _14120_/X _14270_/X vssd1 vssd1 vccd1 vccd1 _18451_/D sky130_fd_sc_hd__o21a_1
X_11483_ _11585_/A vssd1 vssd1 vccd1 vccd1 _14543_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16010_ _14964_/X _19003_/Q _16016_/S vssd1 vssd1 vccd1 vccd1 _16011_/A sky130_fd_sc_hd__mux2_1
XANTENNA_input71_A io_irq_uart_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13222_ _11406_/D _19477_/Q _13222_/S vssd1 vssd1 vccd1 vccd1 _13222_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10434_ _10428_/A _10433_/X _09459_/X vssd1 vssd1 vccd1 vccd1 _10434_/X sky130_fd_sc_hd__o21a_1
XFILLER_171_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12491__B _12495_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13153_ _19826_/Q vssd1 vssd1 vccd1 vccd1 _18119_/B sky130_fd_sc_hd__clkbuf_2
X_10365_ _10365_/A vssd1 vssd1 vccd1 vccd1 _10366_/A sky130_fd_sc_hd__buf_4
XANTENNA__10283__S1 _09486_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10292__A _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _14555_/A _12026_/X _12126_/A _12486_/A vssd1 vssd1 vccd1 vccd1 _12105_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_97_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17961_ _19771_/Q _17963_/C _17960_/Y vssd1 vssd1 vccd1 vccd1 _19771_/D sky130_fd_sc_hd__o21a_1
X_13084_ _19863_/Q _12651_/A _12528_/A _19831_/Q _13083_/X vssd1 vssd1 vccd1 vccd1
+ _13084_/X sky130_fd_sc_hd__a221o_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _18442_/Q vssd1 vssd1 vccd1 vccd1 _10296_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15294__S _15300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14874__A1 _18440_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16912_ _16912_/A vssd1 vssd1 vccd1 vccd1 _19367_/D sky130_fd_sc_hd__clkbuf_1
X_19700_ _19700_/CLK _19700_/D vssd1 vssd1 vccd1 vccd1 _19700_/Q sky130_fd_sc_hd__dfxtp_1
X_12035_ _12035_/A _13607_/A vssd1 vssd1 vccd1 vccd1 _12036_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17892_ _17892_/A vssd1 vssd1 vccd1 vccd1 _17909_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_78_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_124_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19631_ _19631_/CLK _19631_/D vssd1 vssd1 vccd1 vccd1 _19631_/Q sky130_fd_sc_hd__dfxtp_1
X_16843_ _16843_/A vssd1 vssd1 vccd1 vccd1 _19337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19562_ _19626_/CLK _19562_/D vssd1 vssd1 vccd1 vccd1 _19562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16774_ _16774_/A vssd1 vssd1 vccd1 vccd1 _16774_/X sky130_fd_sc_hd__clkbuf_2
X_13986_ _14182_/A _13983_/X _13985_/Y _13894_/A vssd1 vssd1 vccd1 vccd1 _13986_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_65_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13712__C_N _13720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18513_ _18519_/CLK _18513_/D vssd1 vssd1 vccd1 vccd1 _18513_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15725_ _15725_/A vssd1 vssd1 vccd1 vccd1 _18875_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12937_ _18289_/Q _12939_/C _12936_/X vssd1 vssd1 vccd1 vccd1 _18289_/D sky130_fd_sc_hd__a21boi_1
X_19493_ _19786_/CLK _19493_/D vssd1 vssd1 vccd1 vccd1 _19493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12947__A _12983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17014__S _17014_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18444_ _19078_/CLK _18444_/D vssd1 vssd1 vccd1 vccd1 _18444_/Q sky130_fd_sc_hd__dfxtp_4
X_15656_ _18845_/Q _15580_/X _15658_/S vssd1 vssd1 vccd1 vccd1 _15657_/A sky130_fd_sc_hd__mux2_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _18269_/Q _12864_/C _12867_/Y vssd1 vssd1 vccd1 vccd1 _18269_/D sky130_fd_sc_hd__o21a_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15051__A1 _13411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _14513_/A _13106_/B _14603_/X input59/X vssd1 vssd1 vccd1 vccd1 _14608_/B
+ sky130_fd_sc_hd__a22o_1
X_18375_ _19690_/CLK _18375_/D vssd1 vssd1 vccd1 vccd1 _18375_/Q sky130_fd_sc_hd__dfxtp_2
X_11819_ _11706_/X _11816_/X _11818_/X _12696_/A vssd1 vssd1 vccd1 vccd1 _11819_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17328__A0 _16755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15587_ _18815_/Q _15586_/X _15590_/S vssd1 vssd1 vccd1 vccd1 _15588_/A sky130_fd_sc_hd__mux2_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _19872_/Q _19871_/Q _19870_/Q _18242_/A vssd1 vssd1 vccd1 vccd1 _12813_/D
+ sky130_fd_sc_hd__and4_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17326_ _16752_/X _19535_/Q _17330_/S vssd1 vssd1 vccd1 vccd1 _17327_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14538_ _16357_/B _14582_/B vssd1 vssd1 vccd1 vccd1 _14538_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11612__A1 _14553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17257_ _17257_/A vssd1 vssd1 vccd1 vccd1 _19504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14469_ _14469_/A vssd1 vssd1 vccd1 vccd1 _18505_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_49_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_170_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19636_/CLK sky130_fd_sc_hd__clkbuf_16
X_16208_ _16208_/A vssd1 vssd1 vccd1 vccd1 _19076_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17188_ _18440_/Q _13294_/X _17201_/S vssd1 vssd1 vccd1 vccd1 _17188_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16139_ _16213_/B _16920_/B vssd1 vssd1 vccd1 vccd1 _16196_/A sky130_fd_sc_hd__nand2_2
XFILLER_142_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11128__B1 _09625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_185_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19444_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19829_ _19833_/CLK _19829_/D vssd1 vssd1 vccd1 vccd1 _19829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10351__A1 _09171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17713__A _17730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09513_ _10887_/A vssd1 vssd1 vccd1 vccd1 _09514_/A sky130_fd_sc_hd__buf_2
XFILLER_25_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09444_ _11097_/A _09444_/B vssd1 vssd1 vccd1 vccd1 _09444_/X sky130_fd_sc_hd__or2_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_123_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19682_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09231__A _09231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09375_ _11062_/A vssd1 vssd1 vccd1 vccd1 _10950_/A sky130_fd_sc_hd__buf_2
XFILLER_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_138_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19078_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13356__A1 _18292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13356__B2 _18375_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10265__S1 _09697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10150_ _11139_/A _12488_/A vssd1 vssd1 vccd1 vccd1 _11229_/A sky130_fd_sc_hd__or2_1
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10081_ _18773_/Q _19002_/Q _18933_/Q _19231_/Q _09795_/A _10080_/X vssd1 vssd1 vccd1
+ vccd1 _10082_/B sky130_fd_sc_hd__mux4_1
XFILLER_58_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16003__S _16005_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13840_ _13687_/X _13611_/X _13888_/S vssd1 vssd1 vccd1 vccd1 _13840_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15281__A1 _15155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13771_ _13633_/X _13646_/X _13775_/S vssd1 vssd1 vccd1 vccd1 _13771_/X sky130_fd_sc_hd__mux2_1
X_10983_ _18850_/Q _19308_/Q _10983_/S vssd1 vssd1 vccd1 vccd1 _10983_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15510_ _16765_/A vssd1 vssd1 vccd1 vccd1 _15510_/X sky130_fd_sc_hd__clkbuf_2
X_12722_ _19671_/Q _13251_/A _12721_/X vssd1 vssd1 vccd1 vccd1 _12722_/X sky130_fd_sc_hd__a21o_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16490_ _16490_/A vssd1 vssd1 vccd1 vccd1 _19204_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15441_ _15441_/A vssd1 vssd1 vccd1 vccd1 _18763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12653_ _19812_/Q _12518_/A _12602_/A _18323_/Q vssd1 vssd1 vccd1 vccd1 _14946_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18160_ _19840_/Q _18158_/B _18159_/Y vssd1 vssd1 vccd1 vccd1 _19840_/D sky130_fd_sc_hd__o21a_1
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11604_ _13570_/A _13570_/B _13585_/A _13572_/A vssd1 vssd1 vccd1 vccd1 _11604_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15372_ _15372_/A vssd1 vssd1 vccd1 vccd1 _18734_/D sky130_fd_sc_hd__clkbuf_1
X_12584_ _12584_/A vssd1 vssd1 vccd1 vccd1 _12584_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17111_ _16809_/X _19455_/Q _17119_/S vssd1 vssd1 vccd1 vccd1 _17112_/A sky130_fd_sc_hd__mux2_1
X_14323_ _14323_/A _14323_/B vssd1 vssd1 vccd1 vccd1 _14323_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13598__A _13598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18091_ _19816_/Q _18088_/B _18090_/Y vssd1 vssd1 vccd1 vccd1 _19816_/D sky130_fd_sc_hd__o21a_1
X_11535_ _11535_/A vssd1 vssd1 vccd1 vccd1 _12277_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_128_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_50_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17042_ _17042_/A vssd1 vssd1 vccd1 vccd1 _19424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14254_ _14312_/A _14249_/X _14253_/X _13864_/A vssd1 vssd1 vccd1 vccd1 _14254_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_137_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11466_ _15095_/A vssd1 vssd1 vccd1 vccd1 _14173_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_165_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13205_ _13205_/A vssd1 vssd1 vccd1 vccd1 _15242_/D sky130_fd_sc_hd__clkbuf_2
X_10417_ _18598_/Q _19287_/Q _10417_/S vssd1 vssd1 vccd1 vccd1 _10417_/X sky130_fd_sc_hd__mux2_1
X_11397_ _18545_/Q _18544_/Q _18543_/Q _18542_/Q vssd1 vssd1 vccd1 vccd1 _11404_/A
+ sky130_fd_sc_hd__or4b_2
X_14185_ _12142_/A _13933_/A _14184_/X vssd1 vssd1 vccd1 vccd1 _14185_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__16702__A _16702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13136_ _13121_/X _13122_/Y _13134_/X _13135_/X _18619_/Q vssd1 vssd1 vccd1 vccd1
+ _13136_/X sky130_fd_sc_hd__a32o_4
XFILLER_98_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _18600_/Q _19289_/Q _10348_/S vssd1 vssd1 vccd1 vccd1 _10349_/B sky130_fd_sc_hd__mux2_1
XFILLER_97_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18993_ _19414_/CLK _18993_/D vssd1 vssd1 vccd1 vccd1 _18993_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10008__S1 _09147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17944_ _19766_/Q _17944_/B _17944_/C vssd1 vssd1 vccd1 vccd1 _17945_/C sky130_fd_sc_hd__and3_1
X_13067_ _18332_/Q _13067_/B _13067_/C vssd1 vssd1 vccd1 vccd1 _13068_/C sky130_fd_sc_hd__and3_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _18602_/Q _19291_/Q _10279_/S vssd1 vssd1 vccd1 vccd1 _10280_/B sky130_fd_sc_hd__mux2_1
XFILLER_97_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12018_ _11847_/X _12016_/X _12017_/X _11560_/X vssd1 vssd1 vccd1 vccd1 _12018_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09316__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17875_ _17875_/A vssd1 vssd1 vccd1 vccd1 _19738_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17797__A0 _15155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19614_ _19614_/CLK _19614_/D vssd1 vssd1 vccd1 vccd1 _19614_/Q sky130_fd_sc_hd__dfxtp_1
X_16826_ _16826_/A vssd1 vssd1 vccd1 vccd1 _16839_/S sky130_fd_sc_hd__buf_4
XFILLER_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19545_ _19609_/CLK _19545_/D vssd1 vssd1 vccd1 vccd1 _19545_/Q sky130_fd_sc_hd__dfxtp_1
X_16757_ _16757_/A vssd1 vssd1 vccd1 vccd1 _19310_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_40_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19625_/CLK sky130_fd_sc_hd__clkbuf_16
X_13969_ _13968_/X _13814_/Y _13969_/S vssd1 vssd1 vccd1 vccd1 _13969_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15708_ _18868_/Q _15551_/X _15708_/S vssd1 vssd1 vccd1 vccd1 _15709_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11833__A1 _10732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19476_ _19682_/CLK _19476_/D vssd1 vssd1 vccd1 vccd1 _19476_/Q sky130_fd_sc_hd__dfxtp_1
X_16688_ _16688_/A vssd1 vssd1 vccd1 vccd1 _19289_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11833__B2 _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_0_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_15639_ _18837_/Q _15554_/X _15647_/S vssd1 vssd1 vccd1 vccd1 _15640_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18427_ _18818_/CLK _18427_/D vssd1 vssd1 vccd1 vccd1 _18427_/Q sky130_fd_sc_hd__dfxtp_4
X_09160_ _10154_/S vssd1 vssd1 vccd1 vccd1 _10011_/S sky130_fd_sc_hd__clkbuf_4
X_18358_ _18395_/CLK _18358_/D vssd1 vssd1 vccd1 vccd1 _18358_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_55_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19620_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09885__S0 _09866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17309_ _19528_/Q _16728_/X _17313_/S vssd1 vssd1 vccd1 vccd1 _17310_/A sky130_fd_sc_hd__mux2_1
X_09091_ _11585_/B vssd1 vssd1 vccd1 vccd1 _13526_/A sky130_fd_sc_hd__clkbuf_2
X_18289_ _18298_/CLK _18289_/D vssd1 vssd1 vccd1 vccd1 _18289_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__10495__S1 _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13338__A1 _18289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09637__S0 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15927__S _15935_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10247__S1 _09483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11862__A1_N _12473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09993_ _19651_/Q _19068_/Q _19105_/Q _18711_/Q _09983_/X _09763_/A vssd1 vssd1 vccd1
+ vccd1 _09993_/X sky130_fd_sc_hd__mux4_2
XFILLER_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10572__A1 _10475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13510__A1 _13423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15662__S _15662_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12077__A1 _19743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09427_ _09427_/A vssd1 vssd1 vccd1 vccd1 _09428_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16493__S _16497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14774__A0 _14772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09358_ _10329_/A vssd1 vssd1 vccd1 vccd1 _11189_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_139_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09289_ _18577_/Q _18576_/Q _18575_/Q _18574_/Q vssd1 vssd1 vccd1 vccd1 _11665_/B
+ sky130_fd_sc_hd__or4_2
XANTENNA__13211__A _18625_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11320_ _11320_/A vssd1 vssd1 vccd1 vccd1 _14524_/A sky130_fd_sc_hd__inv_2
XFILLER_125_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_2_0_clock clkbuf_4_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_2_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10554__B _10554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15837__S _15841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11251_ _11251_/A vssd1 vssd1 vccd1 vccd1 _11251_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14741__S _14762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10012__B1 _10093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10202_ _09173_/A _10201_/X _09995_/A vssd1 vssd1 vccd1 vccd1 _10202_/X sky130_fd_sc_hd__a21o_1
XFILLER_134_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11182_ _11178_/A _11181_/X _09616_/X vssd1 vssd1 vccd1 vccd1 _11182_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_162_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11666__A _11749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ _10132_/A _10130_/Y _10132_/Y _10177_/A vssd1 vssd1 vccd1 vccd1 _10133_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15138__A _17463_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15990_ _14856_/X _18994_/Q _15994_/S vssd1 vssd1 vccd1 vccd1 _15991_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10064_ _10064_/A _10064_/B vssd1 vssd1 vccd1 vccd1 _10064_/X sky130_fd_sc_hd__or2_1
XANTENNA_input34_A io_ibus_inst[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14941_ _14940_/X _18605_/Q _14941_/S vssd1 vssd1 vccd1 vccd1 _14942_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16668__S _16671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15572__S _15584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17660_ _19669_/Q _17658_/X _17681_/S vssd1 vssd1 vccd1 vccd1 _17661_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09720__A3 _09719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14872_ _17683_/A _14871_/B _14829_/B vssd1 vssd1 vccd1 vccd1 _14872_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16611_ _19261_/Q vssd1 vssd1 vccd1 vccd1 _16612_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__12068__A1 _12043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13823_ _13823_/A vssd1 vssd1 vccd1 vccd1 _13823_/X sky130_fd_sc_hd__clkbuf_2
X_17591_ _17591_/A vssd1 vssd1 vccd1 vccd1 _19653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09469__C1 _09459_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12497__A _12497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19330_ _19331_/CLK _19330_/D vssd1 vssd1 vccd1 vccd1 _19330_/Q sky130_fd_sc_hd__dfxtp_1
X_16542_ _16542_/A vssd1 vssd1 vccd1 vccd1 _19227_/D sky130_fd_sc_hd__clkbuf_1
X_13754_ _13679_/X _13688_/X _13757_/S vssd1 vssd1 vccd1 vccd1 _13754_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10966_ _19246_/Q _19017_/Q _18948_/Q _19342_/Q _10664_/S _10365_/A vssd1 vssd1 vccd1
+ vccd1 _10966_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10174__S0 _10131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12705_ _18278_/Q _12606_/A _12674_/A _18394_/Q _12704_/X vssd1 vssd1 vccd1 vccd1
+ _12705_/X sky130_fd_sc_hd__a221o_1
XANTENNA__17499__S _17507_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19261_ _19616_/CLK _19261_/D vssd1 vssd1 vccd1 vccd1 _19261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16473_ _16093_/X _19197_/Q _16475_/S vssd1 vssd1 vccd1 vccd1 _16474_/A sky130_fd_sc_hd__mux2_1
X_13685_ _14168_/B _14126_/B _13685_/S vssd1 vssd1 vccd1 vccd1 _13685_/X sky130_fd_sc_hd__mux2_1
X_10897_ _10803_/A _10896_/X _10774_/X vssd1 vssd1 vccd1 vccd1 _10897_/Y sky130_fd_sc_hd__o21ai_1
X_18212_ _18223_/A _18212_/B vssd1 vssd1 vccd1 vccd1 _18212_/Y sky130_fd_sc_hd__nor2_1
X_15424_ _18756_/Q _15149_/X _15426_/S vssd1 vssd1 vccd1 vccd1 _15425_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12636_ _13415_/A _18639_/Q vssd1 vssd1 vccd1 vccd1 _12636_/Y sky130_fd_sc_hd__nand2_1
X_19192_ _19709_/CLK _19192_/D vssd1 vssd1 vccd1 vccd1 _19192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18143_ _18159_/A _18148_/C vssd1 vssd1 vccd1 vccd1 _18143_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15355_ _15355_/A vssd1 vssd1 vccd1 vccd1 _18726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12567_ _12567_/A vssd1 vssd1 vccd1 vccd1 _15242_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_129_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16506__A1 _15487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14306_ _18454_/Q _14305_/X _14306_/S vssd1 vssd1 vccd1 vccd1 _14307_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18074_ _18075_/A _18075_/C _18073_/Y vssd1 vssd1 vccd1 vccd1 _19811_/D sky130_fd_sc_hd__o21a_1
X_11518_ _11628_/A _13524_/C _11628_/C _11517_/X vssd1 vssd1 vccd1 vccd1 _11561_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_157_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15286_ _15286_/A vssd1 vssd1 vccd1 vccd1 _18696_/D sky130_fd_sc_hd__clkbuf_1
X_12498_ _12505_/B vssd1 vssd1 vccd1 vccd1 _12503_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15747__S _15747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17025_ _19417_/Q _16686_/X _17025_/S vssd1 vssd1 vccd1 vccd1 _17026_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14237_ _14241_/A _14241_/B vssd1 vssd1 vccd1 vccd1 _14237_/Y sky130_fd_sc_hd__nor2_1
XFILLER_172_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11449_ _11676_/A vssd1 vssd1 vccd1 vccd1 _11720_/B sky130_fd_sc_hd__clkinv_2
XFILLER_153_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16432__A _16488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14168_ _14168_/A _14168_/B vssd1 vssd1 vccd1 vccd1 _14168_/Y sky130_fd_sc_hd__nor2_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _13442_/C _13442_/D _13119_/C vssd1 vssd1 vccd1 vccd1 _13365_/A sky130_fd_sc_hd__and3_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18976_ _19806_/CLK _18976_/D vssd1 vssd1 vccd1 vccd1 _18976_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _14173_/A vssd1 vssd1 vccd1 vccd1 _14099_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17927_ _19761_/Q _19760_/Q _19823_/Q _17927_/D vssd1 vssd1 vccd1 vccd1 _17936_/D
+ sky130_fd_sc_hd__and4_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17858_ _17858_/A vssd1 vssd1 vccd1 vccd1 _19729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16809_ _16809_/A vssd1 vssd1 vccd1 vccd1 _16809_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17789_ _17789_/A vssd1 vssd1 vccd1 vccd1 _19697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19528_ _19624_/CLK _19528_/D vssd1 vssd1 vccd1 vccd1 _19528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19459_ _19557_/CLK _19459_/D vssd1 vssd1 vccd1 vccd1 _19459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09212_ _09212_/A vssd1 vssd1 vccd1 vccd1 _09689_/A sky130_fd_sc_hd__buf_2
XANTENNA__13559__A1 _09094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09143_ _09695_/A vssd1 vssd1 vccd1 vccd1 _09144_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_148_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11742__A0 _10834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10390__A _10390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09976_ _09976_/A _18871_/Q vssd1 vssd1 vccd1 vccd1 _09976_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09950__A3 _09949_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _10928_/A _10820_/B vssd1 vssd1 vccd1 vccd1 _10820_/X sky130_fd_sc_hd__or2_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10751_ _19507_/Q _19121_/Q _19571_/Q _18727_/Q _10669_/A _10670_/X vssd1 vssd1 vccd1
+ vccd1 _10752_/B sky130_fd_sc_hd__mux4_1
XFILLER_13_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13470_ _13470_/A vssd1 vssd1 vccd1 vccd1 _18394_/D sky130_fd_sc_hd__clkbuf_1
X_10682_ _19508_/Q _19122_/Q _19572_/Q _18728_/Q _10860_/S _09139_/A vssd1 vssd1 vccd1
+ vccd1 _10683_/B sky130_fd_sc_hd__mux4_1
XFILLER_71_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12421_ _13702_/A _14310_/B _12399_/B vssd1 vssd1 vccd1 vccd1 _12422_/B sky130_fd_sc_hd__a21o_1
XFILLER_166_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16951__S _16953_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09623__C1 _09403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15140_ _15239_/S vssd1 vssd1 vccd1 vccd1 _15153_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__10233__B1 _10219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12352_ _12353_/A _12372_/A vssd1 vssd1 vccd1 vccd1 _12354_/A sky130_fd_sc_hd__nor2_1
XANTENNA__17161__A1 _13212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11303_ _14900_/A vssd1 vssd1 vccd1 vccd1 _11305_/A sky130_fd_sc_hd__inv_2
X_15071_ _18457_/Q _13435_/B _15071_/S vssd1 vssd1 vccd1 vccd1 _15071_/X sky130_fd_sc_hd__mux2_1
X_12283_ _12284_/A _14253_/A vssd1 vssd1 vccd1 vccd1 _12285_/A sky130_fd_sc_hd__and2_1
XFILLER_135_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14022_ _14285_/A _14026_/A _13797_/A vssd1 vssd1 vccd1 vccd1 _14022_/X sky130_fd_sc_hd__o21a_1
X_11234_ _11234_/A vssd1 vssd1 vccd1 vccd1 _11234_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18830_ _19640_/CLK _18830_/D vssd1 vssd1 vccd1 vccd1 _18830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11165_ _19657_/Q _19074_/Q _19111_/Q _18717_/Q _11153_/X _10306_/X vssd1 vssd1 vccd1
+ vccd1 _11166_/B sky130_fd_sc_hd__mux4_1
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10116_ _18605_/Q _19294_/Q _10153_/S vssd1 vssd1 vccd1 vccd1 _10116_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15973_ _15973_/A vssd1 vssd1 vccd1 vccd1 _18986_/D sky130_fd_sc_hd__clkbuf_1
X_18761_ _19541_/CLK _18761_/D vssd1 vssd1 vccd1 vccd1 _18761_/Q sky130_fd_sc_hd__dfxtp_1
X_11096_ _19514_/Q _19128_/Q _19578_/Q _18734_/Q _10348_/S _09539_/A vssd1 vssd1 vccd1
+ vccd1 _11097_/B sky130_fd_sc_hd__mux4_1
XFILLER_121_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16398__S _16402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10047_ _10140_/A _10047_/B vssd1 vssd1 vccd1 vccd1 _10047_/X sky130_fd_sc_hd__or2_1
X_17712_ _17720_/C _17710_/Y _17711_/X vssd1 vssd1 vccd1 vccd1 _17712_/Y sky130_fd_sc_hd__a21oi_1
X_14924_ _14960_/A vssd1 vssd1 vccd1 vccd1 _14924_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18692_ _19568_/CLK _18692_/D vssd1 vssd1 vccd1 vccd1 _18692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12939__B _18289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17643_ _19666_/Q _17642_/X _17653_/S vssd1 vssd1 vccd1 vccd1 _17644_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14855_ _16680_/A vssd1 vssd1 vccd1 vccd1 _16784_/A sky130_fd_sc_hd__buf_2
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13116__A _14431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13806_ _13806_/A vssd1 vssd1 vccd1 vccd1 _13806_/X sky130_fd_sc_hd__clkbuf_2
X_17574_ _17574_/A vssd1 vssd1 vccd1 vccd1 _19645_/D sky130_fd_sc_hd__clkbuf_1
X_14786_ _14786_/A _18465_/Q _14786_/C vssd1 vssd1 vccd1 vccd1 _14796_/B sky130_fd_sc_hd__and3_1
X_11998_ _11993_/X _11996_/Y _11997_/X vssd1 vssd1 vccd1 vccd1 _11998_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16525_ _19220_/Q _15519_/X _16525_/S vssd1 vssd1 vccd1 vccd1 _16526_/A sky130_fd_sc_hd__mux2_1
X_19313_ _19539_/CLK _19313_/D vssd1 vssd1 vccd1 vccd1 _19313_/Q sky130_fd_sc_hd__dfxtp_1
X_13737_ _13737_/A vssd1 vssd1 vccd1 vccd1 _14054_/A sky130_fd_sc_hd__clkbuf_2
X_10949_ _18820_/Q _19374_/Q _19536_/Q _18788_/Q _10719_/X _09481_/A vssd1 vssd1 vccd1
+ vccd1 _10950_/B sky130_fd_sc_hd__mux4_1
XANTENNA__17924__B1 _19760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09862__C1 _09231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16456_ _16067_/X _19189_/Q _16464_/S vssd1 vssd1 vccd1 vccd1 _16457_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14738__B1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19244_ _19630_/CLK _19244_/D vssd1 vssd1 vccd1 vccd1 _19244_/Q sky130_fd_sc_hd__dfxtp_1
X_13668_ _12381_/A _13667_/X _13668_/S vssd1 vssd1 vccd1 vccd1 _13668_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15407_ _15407_/A vssd1 vssd1 vccd1 vccd1 _18750_/D sky130_fd_sc_hd__clkbuf_1
X_12619_ _13415_/A _18638_/Q vssd1 vssd1 vccd1 vccd1 _12619_/Y sky130_fd_sc_hd__nand2_1
X_19175_ _19724_/CLK _19175_/D vssd1 vssd1 vccd1 vccd1 _19175_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10978__A1_N _18429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16387_ _19159_/Q _15529_/X _16391_/S vssd1 vssd1 vccd1 vccd1 _16388_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10475__A _10475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16861__S _16869_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13599_ _13643_/A vssd1 vssd1 vccd1 vccd1 _13681_/S sky130_fd_sc_hd__buf_2
XFILLER_145_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18126_ _18170_/A vssd1 vssd1 vccd1 vccd1 _18126_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13961__A1 _11787_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15338_ _15338_/A vssd1 vssd1 vccd1 vccd1 _18720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15477__S _15481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18057_ _18059_/A _18059_/C _18039_/X vssd1 vssd1 vccd1 vccd1 _18057_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15269_ _15337_/S vssd1 vssd1 vccd1 vccd1 _15278_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_160_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10870__S1 _10365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17008_ _19409_/Q _16661_/X _17014_/S vssd1 vssd1 vccd1 vccd1 _17009_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11724__B1 _11723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09830_ _09826_/A _09821_/Y _09826_/Y _09942_/A vssd1 vssd1 vccd1 vccd1 _09830_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _09978_/A vssd1 vssd1 vccd1 vccd1 _09984_/A sky130_fd_sc_hd__clkbuf_2
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18959_ _19609_/CLK _18959_/D vssd1 vssd1 vccd1 vccd1 _18959_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16101__S _16113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_172_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09692_ _09692_/A vssd1 vssd1 vccd1 vccd1 _10257_/S sky130_fd_sc_hd__buf_4
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10160__C1 _09230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15940__S _15946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09853__C1 _09231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12204__A1 _12057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10194__A2_N _09309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09126_ _11339_/C vssd1 vssd1 vccd1 vccd1 _11374_/A sky130_fd_sc_hd__buf_2
XANTENNA__17143__A1 _13149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_97_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15387__S _15395_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10518__A1 _09529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09923__A3 _09922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09959_ _18775_/Q _19004_/Q _18935_/Q _19233_/Q _09872_/S _09869_/A vssd1 vssd1 vccd1
+ vccd1 _09960_/B sky130_fd_sc_hd__mux4_1
XFILLER_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14958__C _14958_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ _12972_/A _12972_/B _12969_/Y vssd1 vssd1 vccd1 vccd1 _18304_/D sky130_fd_sc_hd__o21a_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09414__A _09414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ _11922_/A _13614_/A vssd1 vssd1 vccd1 vccd1 _11921_/Y sky130_fd_sc_hd__nand2_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15135__B _16357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10297__A3 _10295_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15850__S _15852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14640_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14640_/X sky130_fd_sc_hd__clkbuf_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _11846_/Y _11851_/Y _12389_/S vssd1 vssd1 vccd1 vccd1 _11852_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _10803_/A _10803_/B vssd1 vssd1 vccd1 vccd1 _10803_/X sky130_fd_sc_hd__or2_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _12533_/A _14564_/X _14570_/Y _14560_/X vssd1 vssd1 vccd1 vccd1 _18545_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12443__A1 _12505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _11783_/A _11783_/B vssd1 vssd1 vccd1 vccd1 _11787_/A sky130_fd_sc_hd__nor2_2
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16310_ _16067_/X _19125_/Q _16318_/S vssd1 vssd1 vccd1 vccd1 _16311_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13522_ _11550_/B _12471_/C _11482_/B vssd1 vssd1 vccd1 vccd1 _13522_/X sky130_fd_sc_hd__o21a_1
X_10734_ _10996_/A vssd1 vssd1 vccd1 vccd1 _10871_/A sky130_fd_sc_hd__clkbuf_2
X_17290_ _17290_/A vssd1 vssd1 vccd1 vccd1 _19519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16241_ _16241_/A vssd1 vssd1 vccd1 vccd1 _19094_/D sky130_fd_sc_hd__clkbuf_1
X_13453_ _18387_/Q _13182_/X _13453_/S vssd1 vssd1 vccd1 vccd1 _13454_/A sky130_fd_sc_hd__mux2_1
X_10665_ _10366_/A _10664_/X _10830_/A vssd1 vssd1 vccd1 vccd1 _10665_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__16681__S _16687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12404_ _12428_/A _12404_/B vssd1 vssd1 vccd1 vccd1 _12406_/A sky130_fd_sc_hd__or2_2
XFILLER_127_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16172_ _16080_/X _19060_/Q _16172_/S vssd1 vssd1 vccd1 vccd1 _16173_/A sky130_fd_sc_hd__mux2_1
X_13384_ _18330_/Q _12663_/X _12665_/A _19819_/Q _13383_/X vssd1 vssd1 vccd1 vccd1
+ _13384_/X sky130_fd_sc_hd__a221o_1
XFILLER_12_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10596_ _10638_/A _10596_/B vssd1 vssd1 vccd1 vccd1 _10596_/X sky130_fd_sc_hd__or2_1
XANTENNA__10301__S0 _09701_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15123_ _15123_/A vssd1 vssd1 vccd1 vccd1 _15123_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12335_ _19753_/Q _19754_/Q _12335_/C vssd1 vssd1 vccd1 vccd1 _12387_/C sky130_fd_sc_hd__and3_1
XFILLER_127_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10852__S1 _09512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11631__A1_N _11997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15054_ _16734_/A vssd1 vssd1 vccd1 vccd1 _16838_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12266_ _12246_/A _12267_/C _19751_/Q vssd1 vssd1 vccd1 vccd1 _12268_/A sky130_fd_sc_hd__a21oi_1
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14214__B _14216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14005_ _14297_/A _14005_/B vssd1 vssd1 vccd1 vccd1 _14005_/X sky130_fd_sc_hd__or2_1
XFILLER_141_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11217_ _13526_/B _11213_/X _11216_/X vssd1 vssd1 vccd1 vccd1 _11217_/X sky130_fd_sc_hd__o21ba_1
X_19862_ _19872_/CLK _19862_/D vssd1 vssd1 vccd1 vccd1 _19862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12197_ _18370_/Q vssd1 vssd1 vccd1 vccd1 _13322_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_122_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12015__A _12043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11182__A1 _11178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15448__A1 _15184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput81 _12115_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[17] sky130_fd_sc_hd__buf_2
XFILLER_95_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18813_ _19657_/CLK _18813_/D vssd1 vssd1 vccd1 vccd1 _18813_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput92 _12358_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[27] sky130_fd_sc_hd__buf_2
XFILLER_95_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11148_ _11148_/A _12497_/A vssd1 vssd1 vccd1 vccd1 _11149_/B sky130_fd_sc_hd__nor2_1
XFILLER_96_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19793_ _19795_/CLK _19793_/D vssd1 vssd1 vccd1 vccd1 _19793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17017__S _17025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18744_ _19427_/CLK _18744_/D vssd1 vssd1 vccd1 vccd1 _18744_/Q sky130_fd_sc_hd__dfxtp_1
X_11079_ _11248_/A _11248_/B _11248_/C vssd1 vssd1 vccd1 vccd1 _11080_/C sky130_fd_sc_hd__a21o_1
X_15956_ _17779_/A _15956_/B vssd1 vssd1 vccd1 vccd1 _15957_/A sky130_fd_sc_hd__and2_2
XFILLER_36_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14907_ _16693_/A vssd1 vssd1 vccd1 vccd1 _16797_/A sky130_fd_sc_hd__clkbuf_2
X_18675_ _19720_/CLK _18675_/D vssd1 vssd1 vccd1 vccd1 _18675_/Q sky130_fd_sc_hd__dfxtp_1
X_15887_ _14740_/X _18947_/Q _15891_/S vssd1 vssd1 vccd1 vccd1 _15888_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17626_ _17626_/A vssd1 vssd1 vccd1 vccd1 _19663_/D sky130_fd_sc_hd__clkbuf_1
X_14838_ _14838_/A vssd1 vssd1 vccd1 vccd1 _14838_/X sky130_fd_sc_hd__buf_2
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17557_ _19638_/Q _16774_/A _17557_/S vssd1 vssd1 vccd1 vccd1 _17558_/A sky130_fd_sc_hd__mux2_1
X_14769_ _14766_/Y _14768_/X _14923_/S vssd1 vssd1 vccd1 vccd1 _14769_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16508_ _19212_/Q _15494_/X _16514_/S vssd1 vssd1 vccd1 vccd1 _16509_/A sky130_fd_sc_hd__mux2_1
X_17488_ _19607_/Q _16673_/X _17496_/S vssd1 vssd1 vccd1 vccd1 _17489_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19227_ _19642_/CLK _19227_/D vssd1 vssd1 vccd1 vccd1 _19227_/Q sky130_fd_sc_hd__dfxtp_1
X_16439_ _16439_/A vssd1 vssd1 vccd1 vccd1 _19181_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10409__S _10494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_119_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13934__A1 _11751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19158_ _19707_/CLK _19158_/D vssd1 vssd1 vccd1 vccd1 _19158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18109_ _18110_/B _18110_/C _19824_/Q vssd1 vssd1 vccd1 vccd1 _18111_/B sky130_fd_sc_hd__a21oi_1
XFILLER_117_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10843__S1 _10785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19089_ _19635_/CLK _19089_/D vssd1 vssd1 vccd1 vccd1 _19089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14124__B _14126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15935__S _15935_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11173__A1 _09689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09813_ _18841_/Q _19395_/Q _19557_/Q _18809_/Q _09928_/A _09875_/A vssd1 vssd1 vccd1
+ vccd1 _09814_/B sky130_fd_sc_hd__mux4_1
XFILLER_141_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09744_ _19655_/Q _19072_/Q _19109_/Q _18715_/Q _09721_/X _09723_/X vssd1 vssd1 vccd1
+ vccd1 _09744_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09675_ _18613_/Q _19302_/Q _09675_/S vssd1 vssd1 vccd1 vccd1 _09676_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10133__C1 _10177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12595__A _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17597__S _17601_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10450_ _18598_/Q _19287_/Q _10450_/S vssd1 vssd1 vccd1 vccd1 _10451_/B sky130_fd_sc_hd__mux2_1
XFILLER_164_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09109_ _11528_/A _09113_/A vssd1 vssd1 vccd1 vccd1 _09109_/Y sky130_fd_sc_hd__nor2_4
X_10381_ _09640_/A _10380_/X _09708_/A vssd1 vssd1 vccd1 vccd1 _10381_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10601__A_N _12474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15678__A1 _15506_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12120_ _19676_/Q _11563_/X _11560_/X vssd1 vssd1 vccd1 vccd1 _12120_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09409__A _09409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13689__A0 _14176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12051_ _13295_/A _12075_/C vssd1 vssd1 vccd1 vccd1 _12051_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11164__A1 _09689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11002_ _18850_/Q _19308_/Q _11051_/S vssd1 vssd1 vccd1 vccd1 _11003_/B sky130_fd_sc_hd__mux2_1
XFILLER_89_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10372__C1 _09459_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15810_ _15878_/S vssd1 vssd1 vccd1 vccd1 _15819_/S sky130_fd_sc_hd__clkbuf_4
X_16790_ _16790_/A vssd1 vssd1 vccd1 vccd1 _16790_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12376__A1_N _11517_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13310__C1 _13282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12489__B _12495_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15741_ _14729_/X _18882_/Q _15747_/S vssd1 vssd1 vccd1 vccd1 _15742_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09144__A _09144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ _12983_/A _12953_/B _12957_/C vssd1 vssd1 vccd1 vccd1 _18294_/D sky130_fd_sc_hd__nor3_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14985__A _16715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ _19668_/Q _11959_/B vssd1 vssd1 vccd1 vccd1 _11904_/X sky130_fd_sc_hd__or2_1
XFILLER_46_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15672_ _15672_/A vssd1 vssd1 vccd1 vccd1 _18851_/D sky130_fd_sc_hd__clkbuf_1
X_18460_ _18623_/CLK _18460_/D vssd1 vssd1 vccd1 vccd1 _18460_/Q sky130_fd_sc_hd__dfxtp_1
X_12884_ _12904_/A _12884_/B _12884_/C vssd1 vssd1 vccd1 vccd1 _18274_/D sky130_fd_sc_hd__nor3_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _18562_/Q _14613_/X _14622_/X input64/X vssd1 vssd1 vccd1 vccd1 _14624_/B
+ sky130_fd_sc_hd__a22o_1
X_17411_ _16771_/X _19573_/Q _17413_/S vssd1 vssd1 vccd1 vccd1 _17412_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18391_ _19690_/CLK _18391_/D vssd1 vssd1 vccd1 vccd1 _18391_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _11834_/X _11738_/A _11835_/S vssd1 vssd1 vccd1 vccd1 _13761_/A sky130_fd_sc_hd__mux2_2
XANTENNA__09817__C1 _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17342_/A vssd1 vssd1 vccd1 vccd1 _19542_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _18538_/Q _14550_/X _14553_/X _14548_/X vssd1 vssd1 vccd1 vccd1 _18538_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _18354_/Q _15255_/A vssd1 vssd1 vccd1 vccd1 _11766_/X sky130_fd_sc_hd__or2_1
XFILLER_159_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13505_ _13505_/A vssd1 vssd1 vccd1 vccd1 _18410_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17273_ _17273_/A vssd1 vssd1 vccd1 vccd1 _19511_/D sky130_fd_sc_hd__clkbuf_1
X_10717_ _11056_/A vssd1 vssd1 vccd1 vccd1 _10807_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14485_ _18513_/Q _19751_/Q _14487_/S vssd1 vssd1 vccd1 vccd1 _14486_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_120_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11697_ _11696_/Y _18493_/Q _11697_/S vssd1 vssd1 vccd1 vccd1 _13667_/A sky130_fd_sc_hd__mux2_4
XFILLER_158_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16705__A _16705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17300__S _17302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16224_ _16048_/X _19087_/Q _16224_/S vssd1 vssd1 vccd1 vccd1 _16225_/A sky130_fd_sc_hd__mux2_1
X_19012_ _19285_/CLK _19012_/D vssd1 vssd1 vccd1 vccd1 _19012_/Q sky130_fd_sc_hd__dfxtp_1
X_13436_ _12556_/X _13426_/Y _13435_/X _12712_/X _18650_/Q vssd1 vssd1 vccd1 vccd1
+ _15262_/B sky130_fd_sc_hd__a32oi_4
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10648_ _18857_/Q _19315_/Q _10648_/S vssd1 vssd1 vccd1 vccd1 _10649_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12952__B _18293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11849__A _11849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16155_ _16055_/X _19052_/Q _16161_/S vssd1 vssd1 vccd1 vccd1 _16156_/A sky130_fd_sc_hd__mux2_1
X_13367_ _13354_/X _13364_/X _13366_/X _13350_/X vssd1 vssd1 vccd1 vccd1 _18375_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10579_ _18858_/Q _19316_/Q _10579_/S vssd1 vssd1 vccd1 vccd1 _10580_/B sky130_fd_sc_hd__mux2_1
XFILLER_155_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15669__A1 _15494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15106_ _18630_/Q _15102_/X _15104_/X _11082_/B vssd1 vssd1 vccd1 vccd1 _18630_/D
+ sky130_fd_sc_hd__a22o_1
X_12318_ _11980_/X _12316_/X _12317_/X vssd1 vssd1 vccd1 vccd1 _12318_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_154_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16086_ _16086_/A vssd1 vssd1 vccd1 vccd1 _19029_/D sky130_fd_sc_hd__clkbuf_1
X_13298_ _13403_/A _18634_/Q vssd1 vssd1 vccd1 vccd1 _13298_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15037_ _18485_/Q _18486_/Q _15037_/C vssd1 vssd1 vccd1 vccd1 _15049_/B sky130_fd_sc_hd__and3_1
X_12249_ _12244_/X _12247_/X _12248_/X _12072_/X vssd1 vssd1 vccd1 vccd1 _12249_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17536__A _17592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19845_ _19866_/CLK _19845_/D vssd1 vssd1 vccd1 vccd1 _19845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19776_ _19858_/CLK _19776_/D vssd1 vssd1 vccd1 vccd1 _19776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16988_ _16841_/X _19401_/Q _16990_/S vssd1 vssd1 vccd1 vccd1 _16989_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_45_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18727_ _19571_/CLK _18727_/D vssd1 vssd1 vccd1 vccd1 _18727_/Q sky130_fd_sc_hd__dfxtp_1
X_15939_ _15939_/A vssd1 vssd1 vccd1 vccd1 _18970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17271__A _17317_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ _09463_/A _09455_/X _09458_/X _09459_/X vssd1 vssd1 vccd1 vccd1 _09460_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18658_ _19442_/CLK _18658_/D vssd1 vssd1 vccd1 vccd1 _18658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10761__S0 _10836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17609_ _17621_/C _17609_/B vssd1 vssd1 vccd1 vccd1 _17609_/Y sky130_fd_sc_hd__nand2_2
X_09391_ _09391_/A vssd1 vssd1 vccd1 vccd1 _09392_/A sky130_fd_sc_hd__clkbuf_4
X_18589_ _19599_/CLK _18589_/D vssd1 vssd1 vccd1 vccd1 _18589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10816__S1 _10969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09229__A _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10004__A_N _10003_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16085__A1 _19029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11494__A _18561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09727_ _09727_/A vssd1 vssd1 vccd1 vccd1 _09727_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12646__A1 _18343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12646__B2 _19489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09658_ _19624_/Q _19462_/Q _18908_/Q _18678_/Q _09342_/A _09603_/A vssd1 vssd1 vccd1
+ vccd1 _09659_/B sky130_fd_sc_hd__mux4_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09589_ _09735_/A vssd1 vssd1 vccd1 vccd1 _09728_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _11619_/Y _18491_/Q _11697_/S vssd1 vssd1 vccd1 vccd1 _13671_/A sky130_fd_sc_hd__mux2_4
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11551_ _11551_/A _11551_/B vssd1 vssd1 vccd1 vccd1 _11551_/Y sky130_fd_sc_hd__nand2_1
XFILLER_168_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10502_ _19608_/Q _19446_/Q _18892_/Q _18662_/Q _10500_/X _10501_/X vssd1 vssd1 vccd1
+ vccd1 _10503_/B sky130_fd_sc_hd__mux4_2
XFILLER_168_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14270_ _12313_/Y _13730_/X _14269_/X _14099_/X vssd1 vssd1 vccd1 vccd1 _14270_/X
+ sky130_fd_sc_hd__a211o_1
X_11482_ _11366_/A _11482_/B _11538_/A _13520_/B vssd1 vssd1 vccd1 vccd1 _11522_/A
+ sky130_fd_sc_hd__and4b_1
X_13221_ _19667_/Q _12624_/A _12742_/A _18391_/Q vssd1 vssd1 vccd1 vccd1 _13221_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10433_ _19609_/Q _19447_/Q _18893_/Q _18663_/Q _09632_/A _10368_/X vssd1 vssd1 vccd1
+ vccd1 _10433_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12491__C _12491_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input64_A io_ibus_inst[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13152_ _13426_/A _18621_/Q vssd1 vssd1 vccd1 vccd1 _13152_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09139__A _09139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10364_ _10364_/A vssd1 vssd1 vccd1 vccd1 _10365_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ _12095_/A _12002_/X _12102_/X vssd1 vssd1 vccd1 vccd1 _12103_/X sky130_fd_sc_hd__o21a_1
XANTENNA__15575__S _15584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17960_ _19771_/Q _17963_/C _17950_/X vssd1 vssd1 vccd1 vccd1 _17960_/Y sky130_fd_sc_hd__a21oi_1
X_13083_ _13078_/X _13079_/X _13082_/X _12628_/A _19767_/Q vssd1 vssd1 vccd1 vccd1
+ _13083_/X sky130_fd_sc_hd__o32a_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10295_ _10288_/Y _10290_/Y _10292_/Y _10294_/Y _09402_/A vssd1 vssd1 vccd1 vccd1
+ _10295_/X sky130_fd_sc_hd__o221a_2
XFILLER_151_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12334__B1 _19754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13531__C1 _13530_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16911_ _19367_/Q _16731_/X _16913_/S vssd1 vssd1 vccd1 vccd1 _16912_/A sky130_fd_sc_hd__mux2_1
X_12034_ _12035_/A _13607_/A vssd1 vssd1 vccd1 vccd1 _12036_/A sky130_fd_sc_hd__and2_1
XFILLER_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17891_ _17891_/A vssd1 vssd1 vccd1 vccd1 _19746_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17790__S _17794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19630_ _19630_/CLK _19630_/D vssd1 vssd1 vccd1 vccd1 _19630_/Q sky130_fd_sc_hd__dfxtp_1
X_16842_ _16841_/X _19337_/Q _16845_/S vssd1 vssd1 vccd1 vccd1 _16843_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10991__S0 _10668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13108__B _13108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19561_ _19657_/CLK _19561_/D vssd1 vssd1 vccd1 vccd1 _19561_/Q sky130_fd_sc_hd__dfxtp_1
X_16773_ _16773_/A vssd1 vssd1 vccd1 vccd1 _19315_/D sky130_fd_sc_hd__clkbuf_1
X_13985_ _14078_/A _13976_/Y _13984_/Y vssd1 vssd1 vccd1 vccd1 _13985_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14919__S _14941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18512_ _18519_/CLK _18512_/D vssd1 vssd1 vccd1 vccd1 _18512_/Q sky130_fd_sc_hd__dfxtp_1
X_12936_ _18289_/Q _12939_/C _17895_/A vssd1 vssd1 vccd1 vccd1 _12936_/X sky130_fd_sc_hd__o21a_1
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15724_ _18875_/Q _15574_/X _15730_/S vssd1 vssd1 vccd1 vccd1 _15725_/A sky130_fd_sc_hd__mux2_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19492_ _19786_/CLK _19492_/D vssd1 vssd1 vccd1 vccd1 _19492_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09602__A _09602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18443_ _19078_/CLK _18443_/D vssd1 vssd1 vccd1 vccd1 _18443_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12867_ _12897_/A _12873_/C vssd1 vssd1 vccd1 vccd1 _12867_/Y sky130_fd_sc_hd__nor2_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15655_ _15655_/A vssd1 vssd1 vccd1 vccd1 _18844_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _19665_/Q _11959_/B vssd1 vssd1 vccd1 vccd1 _11818_/X sky130_fd_sc_hd__or2_1
X_14606_ _14606_/A vssd1 vssd1 vccd1 vccd1 _18556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18374_ _18381_/CLK _18374_/D vssd1 vssd1 vccd1 vccd1 _18374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15586_ _16841_/A vssd1 vssd1 vccd1 vccd1 _15586_/X sky130_fd_sc_hd__clkbuf_2
X_12798_ _19869_/Q _19868_/Q _19867_/Q _18234_/A vssd1 vssd1 vccd1 vccd1 _18242_/A
+ sky130_fd_sc_hd__and4_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14537_ _15412_/B vssd1 vssd1 vccd1 vccd1 _16357_/B sky130_fd_sc_hd__clkbuf_4
X_17325_ _17325_/A vssd1 vssd1 vccd1 vccd1 _19534_/D sky130_fd_sc_hd__clkbuf_1
X_11749_ _11749_/A vssd1 vssd1 vccd1 vccd1 _12016_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17030__S _17036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17256_ _19504_/Q _16651_/X _17258_/S vssd1 vssd1 vccd1 vccd1 _17257_/A sky130_fd_sc_hd__mux2_1
X_14468_ _18505_/Q _19743_/Q _14476_/S vssd1 vssd1 vccd1 vccd1 _14469_/A sky130_fd_sc_hd__mux2_1
X_13419_ _19790_/Q _12629_/S _13417_/X _13418_/X vssd1 vssd1 vccd1 vccd1 _13419_/X
+ sky130_fd_sc_hd__o22a_1
X_16207_ _16131_/X _19076_/Q _16209_/S vssd1 vssd1 vccd1 vccd1 _16208_/A sky130_fd_sc_hd__mux2_1
X_17187_ _17204_/A vssd1 vssd1 vccd1 vccd1 _17201_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_143_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14399_ _17716_/A _18510_/Q _14410_/S vssd1 vssd1 vccd1 vccd1 _14400_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16138_ _16138_/A _16138_/B _16212_/C _16212_/D vssd1 vssd1 vccd1 vccd1 _16920_/B
+ sky130_fd_sc_hd__and4_4
XFILLER_6_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15485__S _15485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16069_ _16067_/X _19024_/Q _16081_/S vssd1 vssd1 vccd1 vccd1 _16070_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11128__A1 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09416__S1 _09364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09741__A1 _09318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19828_ _19833_/CLK _19828_/D vssd1 vssd1 vccd1 vccd1 _19828_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_84_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19759_ _19759_/CLK _19759_/D vssd1 vssd1 vccd1 vccd1 _19759_/Q sky130_fd_sc_hd__dfxtp_4
X_09512_ _09512_/A vssd1 vssd1 vccd1 vccd1 _10887_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09512__A _09512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09443_ _19273_/Q _19044_/Q _18975_/Q _19369_/Q _10350_/S _09442_/X vssd1 vssd1 vccd1
+ vccd1 _09444_/B sky130_fd_sc_hd__mux4_1
XFILLER_80_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13034__A _13034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09374_ _10695_/A vssd1 vssd1 vccd1 vccd1 _11062_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15750__A0 _14772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13210__D1 _13209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15395__S _15395_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14305__A1 _12385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12316__A0 _12313_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16080__A _16790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10080_ _10080_/A vssd1 vssd1 vccd1 vccd1 _10080_/X sky130_fd_sc_hd__buf_4
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17115__S _17119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13770_ _13766_/X _13769_/X _13991_/S vssd1 vssd1 vccd1 vccd1 _13770_/X sky130_fd_sc_hd__mux2_1
X_10982_ _18587_/Q _19276_/Q _10982_/S vssd1 vssd1 vccd1 vccd1 _10982_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12721_ _18395_/Q _12742_/A _12719_/X _12720_/X vssd1 vssd1 vccd1 vccd1 _12721_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_167_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15440_ _18763_/Q _15171_/X _15448_/S vssd1 vssd1 vccd1 vccd1 _15441_/A sky130_fd_sc_hd__mux2_1
X_12652_ _12821_/B _12651_/X _12528_/X _19844_/Q vssd1 vssd1 vccd1 vccd1 _14946_/C
+ sky130_fd_sc_hd__a22o_2
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11603_ _11310_/X _09119_/B _11474_/A vssd1 vssd1 vccd1 vccd1 _13572_/A sky130_fd_sc_hd__a21o_1
XFILLER_30_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15371_ _18734_/Q _15181_/X _15373_/S vssd1 vssd1 vccd1 vccd1 _15372_/A sky130_fd_sc_hd__mux2_1
X_12583_ _12583_/A vssd1 vssd1 vccd1 vccd1 _12584_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12783__A _18533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17110_ _17121_/A vssd1 vssd1 vccd1 vccd1 _17119_/S sky130_fd_sc_hd__buf_4
X_14322_ _14324_/A _14324_/B vssd1 vssd1 vccd1 vccd1 _14323_/B sky130_fd_sc_hd__and2_1
X_18090_ _18114_/A _18094_/C vssd1 vssd1 vccd1 vccd1 _18090_/Y sky130_fd_sc_hd__nor2_1
X_11534_ _11534_/A _11534_/B _11468_/B vssd1 vssd1 vccd1 vccd1 _11535_/A sky130_fd_sc_hd__or3b_4
XFILLER_157_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17041_ _19424_/Q _16709_/X _17047_/S vssd1 vssd1 vccd1 vccd1 _17042_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15741__A0 _14729_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14253_ _14253_/A _12280_/A vssd1 vssd1 vccd1 vccd1 _14253_/X sky130_fd_sc_hd__or2b_1
X_11465_ _14601_/A _13442_/C vssd1 vssd1 vccd1 vccd1 _15095_/A sky130_fd_sc_hd__nand2_2
X_13204_ _12883_/B _12638_/X _13119_/C _18356_/Q vssd1 vssd1 vccd1 vccd1 _13204_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10416_ _10428_/A _10416_/B vssd1 vssd1 vccd1 vccd1 _10416_/X sky130_fd_sc_hd__or2_1
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14184_ _13931_/A _14106_/X _14183_/X _13871_/X vssd1 vssd1 vccd1 vccd1 _14184_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_174_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11396_ _11412_/A _11400_/A _11413_/A vssd1 vssd1 vccd1 vccd1 _13130_/A sky130_fd_sc_hd__nor3_4
XFILLER_48_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13135_ _13306_/A vssd1 vssd1 vccd1 vccd1 _13135_/X sky130_fd_sc_hd__buf_2
XFILLER_174_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10347_ _11135_/A _12483_/A vssd1 vssd1 vccd1 vccd1 _11239_/A sky130_fd_sc_hd__or2_1
XFILLER_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18992_ _19707_/CLK _18992_/D vssd1 vssd1 vccd1 vccd1 _18992_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _17944_/B _17944_/C _19766_/Q vssd1 vssd1 vccd1 vccd1 _17945_/B sky130_fd_sc_hd__a21oi_1
X_13066_ _13067_/B _13067_/C _18332_/Q vssd1 vssd1 vccd1 vccd1 _13068_/B sky130_fd_sc_hd__a21oi_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10278_ _10278_/A vssd1 vssd1 vccd1 vccd1 _10278_/Y sky130_fd_sc_hd__inv_2
X_12017_ _19672_/Q _12017_/B vssd1 vssd1 vccd1 vccd1 _12017_/X sky130_fd_sc_hd__or2_1
XFILLER_94_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10869__B1 _09244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10242__S _10242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17874_ _17874_/A _17874_/B vssd1 vssd1 vccd1 vccd1 _17875_/A sky130_fd_sc_hd__or2_1
XANTENNA__12023__A _14589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19613_ _19613_/CLK _19613_/D vssd1 vssd1 vccd1 vccd1 _19613_/Q sky130_fd_sc_hd__dfxtp_1
X_16825_ _16825_/A vssd1 vssd1 vccd1 vccd1 _16825_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12958__A _12983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17025__S _17025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19544_ _19608_/CLK _19544_/D vssd1 vssd1 vccd1 vccd1 _19544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16756_ _16755_/X _19310_/Q _16759_/S vssd1 vssd1 vccd1 vccd1 _16757_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13968_ _13843_/X _13848_/A _13968_/S vssd1 vssd1 vccd1 vccd1 _13968_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15707_ _15707_/A vssd1 vssd1 vccd1 vccd1 _18867_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12919_ _18284_/Q _12925_/C _12919_/C vssd1 vssd1 vccd1 vccd1 _12930_/D sky130_fd_sc_hd__and3_1
X_19475_ _19689_/CLK _19475_/D vssd1 vssd1 vccd1 vccd1 _19475_/Q sky130_fd_sc_hd__dfxtp_1
X_13899_ _13899_/A vssd1 vssd1 vccd1 vccd1 _13899_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16687_ _19289_/Q _16686_/X _16687_/S vssd1 vssd1 vccd1 vccd1 _16688_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18426_ _19468_/CLK _18426_/D vssd1 vssd1 vccd1 vccd1 _18426_/Q sky130_fd_sc_hd__dfxtp_1
X_15638_ _15649_/A vssd1 vssd1 vccd1 vccd1 _15647_/S sky130_fd_sc_hd__buf_4
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18357_ _18357_/CLK _18357_/D vssd1 vssd1 vccd1 vccd1 _18357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15569_ _15569_/A vssd1 vssd1 vccd1 vccd1 _18809_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09885__S1 _09869_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17308_ _17308_/A vssd1 vssd1 vccd1 vccd1 _19527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09090_ _11376_/C vssd1 vssd1 vccd1 vccd1 _11585_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18288_ _18298_/CLK _18288_/D vssd1 vssd1 vccd1 vccd1 _18288_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_147_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17239_ _19498_/Q hold4/X _17239_/S vssd1 vssd1 vccd1 vccd1 _17240_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10417__S _10417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09992_ _09992_/A _09992_/B vssd1 vssd1 vccd1 vccd1 _09992_/X sky130_fd_sc_hd__or2_1
XANTENNA__16104__S _16113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10660__B _12473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10955__S0 _10909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12077__A2 _11788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09242__A _19695_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11824__A2 _11822_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09426_ _09624_/A _09624_/B _09425_/Y vssd1 vssd1 vccd1 vccd1 _09427_/A sky130_fd_sc_hd__a21o_2
XFILLER_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09357_ _11113_/A vssd1 vssd1 vccd1 vccd1 _10329_/A sky130_fd_sc_hd__buf_2
XFILLER_166_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09288_ _18533_/Q vssd1 vssd1 vccd1 vccd1 _15339_/A sky130_fd_sc_hd__inv_2
XFILLER_138_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_167_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13211__B _13211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12108__A _14168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11250_ _11220_/A _11198_/Y _11249_/Y _09755_/A vssd1 vssd1 vccd1 vccd1 _11250_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_134_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10012__A1 _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10201_ _18866_/Q _19324_/Q _10256_/S vssd1 vssd1 vccd1 vccd1 _10201_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09953__A1 _09810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11181_ _19657_/Q _19074_/Q _19111_/Q _18717_/Q _10185_/S _09736_/A vssd1 vssd1 vccd1
+ vccd1 _11181_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16014__S _16016_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10132_ _10132_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _10132_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16949__S _16953_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10063_ _19521_/Q _19135_/Q _19585_/Q _18741_/Q _09808_/A _09936_/A vssd1 vssd1 vccd1
+ vccd1 _10064_/B sky130_fd_sc_hd__mux4_1
X_14940_ _16806_/A vssd1 vssd1 vccd1 vccd1 _14940_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input27_A io_dbus_rdata[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14871_ _18472_/Q _14871_/B vssd1 vssd1 vccd1 vccd1 _14894_/C sky130_fd_sc_hd__and2_1
XFILLER_85_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16451__A1 _19187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16610_ _16610_/A vssd1 vssd1 vccd1 vccd1 _19260_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13822_ _13893_/A vssd1 vssd1 vccd1 vccd1 _13823_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17590_ _19653_/Q _16822_/A _17590_/S vssd1 vssd1 vccd1 vccd1 _17591_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12068__A2 _12067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09152__A _09152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13753_ _14103_/A vssd1 vssd1 vccd1 vccd1 _13753_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16541_ _19227_/Q _15542_/X _16547_/S vssd1 vssd1 vccd1 vccd1 _16542_/A sky130_fd_sc_hd__mux2_1
X_10965_ _09208_/A _10956_/Y _10958_/Y _10962_/Y _10964_/Y vssd1 vssd1 vccd1 vccd1
+ _10965_/X sky130_fd_sc_hd__o32a_1
XFILLER_43_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16684__S _16687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__A _10299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17400__A0 _16755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10174__S1 _09610_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12704_ _12545_/A _18361_/Q _15242_/B _12640_/A vssd1 vssd1 vccd1 vccd1 _12704_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_43_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19260_ _19613_/CLK _19260_/D vssd1 vssd1 vccd1 vccd1 _19260_/Q sky130_fd_sc_hd__dfxtp_1
X_13684_ _13680_/X _13683_/X _13776_/S vssd1 vssd1 vccd1 vccd1 _13684_/X sky130_fd_sc_hd__mux2_1
X_16472_ _16472_/A vssd1 vssd1 vccd1 vccd1 _19196_/D sky130_fd_sc_hd__clkbuf_1
X_10896_ _19631_/Q _19048_/Q _19085_/Q _18691_/Q _10631_/A _10726_/X vssd1 vssd1 vccd1
+ vccd1 _10896_/X sky130_fd_sc_hd__mux4_2
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18211_ _18214_/B _18214_/C vssd1 vssd1 vccd1 vccd1 _18212_/B sky130_fd_sc_hd__and2_1
X_12635_ _18337_/Q _12574_/X _12575_/X _12634_/X vssd1 vssd1 vccd1 vccd1 _18337_/D
+ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_184_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19706_/CLK sky130_fd_sc_hd__clkbuf_16
X_15423_ _15423_/A vssd1 vssd1 vccd1 vccd1 _18755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19191_ _19609_/CLK _19191_/D vssd1 vssd1 vccd1 vccd1 _19191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18142_ _19834_/Q _19833_/Q _19832_/Q _18142_/D vssd1 vssd1 vccd1 vccd1 _18148_/C
+ sky130_fd_sc_hd__and4_1
X_15354_ _18726_/Q _15155_/X _15362_/S vssd1 vssd1 vccd1 vccd1 _15355_/A sky130_fd_sc_hd__mux2_1
X_12566_ _12566_/A vssd1 vssd1 vccd1 vccd1 _14562_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_129_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10251__A1 _09402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14305_ _12385_/X _14102_/A _14303_/X _14304_/Y vssd1 vssd1 vccd1 vccd1 _14305_/X
+ sky130_fd_sc_hd__a22o_2
X_11517_ _14584_/A _11517_/B _14566_/A _13524_/B vssd1 vssd1 vccd1 vccd1 _11517_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_144_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18073_ _18075_/A _18075_/C _18039_/X vssd1 vssd1 vccd1 vccd1 _18073_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_129_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15285_ _18696_/Q _15162_/X _15289_/S vssd1 vssd1 vccd1 vccd1 _15286_/A sky130_fd_sc_hd__mux2_1
X_12497_ _12497_/A _12497_/B vssd1 vssd1 vccd1 vccd1 _12497_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output95_A _11667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17024_ _17024_/A vssd1 vssd1 vccd1 vccd1 _19416_/D sky130_fd_sc_hd__clkbuf_1
X_14236_ _14236_/A vssd1 vssd1 vccd1 vccd1 _18448_/D sky130_fd_sc_hd__clkbuf_1
X_11448_ _11444_/X _11721_/A _11447_/X _18335_/Q vssd1 vssd1 vccd1 vccd1 _11676_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_144_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14167_ _13927_/X _14164_/Y _14166_/X _13862_/A vssd1 vssd1 vccd1 vccd1 _14167_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_124_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11379_ _11371_/Y _11610_/A _09624_/B vssd1 vssd1 vccd1 vccd1 _11379_/X sky130_fd_sc_hd__a21bo_1
XFILLER_112_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09686__A2_N _09309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13118_ _13311_/A vssd1 vssd1 vccd1 vccd1 _13118_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_122_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19488_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09327__A _10496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14098_ _14054_/X _14086_/X _14096_/X _14097_/X vssd1 vssd1 vccd1 vccd1 _14098_/X
+ sky130_fd_sc_hd__o211a_1
X_18975_ _19550_/CLK _18975_/D vssd1 vssd1 vccd1 vccd1 _18975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15763__S _15769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ _17935_/A _17926_/B _17926_/C vssd1 vssd1 vccd1 vccd1 _19760_/D sky130_fd_sc_hd__nor3_1
X_13049_ _13049_/A _13055_/C vssd1 vssd1 vccd1 vccd1 _13049_/Y sky130_fd_sc_hd__nor2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17857_ _17890_/A _17857_/B vssd1 vssd1 vccd1 vccd1 _17858_/A sky130_fd_sc_hd__and2_1
XFILLER_67_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16808_ _16808_/A vssd1 vssd1 vccd1 vccd1 _19326_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_137_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _18818_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17788_ _15143_/X _19697_/Q _17794_/S vssd1 vssd1 vccd1 vccd1 _17789_/A sky130_fd_sc_hd__mux2_1
X_19527_ _19591_/CLK _19527_/D vssd1 vssd1 vccd1 vccd1 _19527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16739_ _16739_/A vssd1 vssd1 vccd1 vccd1 _19305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19458_ _19556_/CLK _19458_/D vssd1 vssd1 vccd1 vccd1 _19458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09211_ _09434_/A vssd1 vssd1 vccd1 vccd1 _09212_/A sky130_fd_sc_hd__buf_2
XFILLER_61_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18409_ _19689_/CLK _18409_/D vssd1 vssd1 vccd1 vccd1 _18409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19389_ _19715_/CLK _19389_/D vssd1 vssd1 vccd1 vccd1 _19389_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11114__S0 _11110_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09142_ _09142_/A vssd1 vssd1 vccd1 vccd1 _09695_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15938__S _15946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11990__A1 _19671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09396__C1 _09395_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09237__A _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09975_ _09783_/A _09974_/X _10107_/A vssd1 vssd1 vccd1 vccd1 _09975_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13495__A1 _12757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17630__A0 _19664_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12110__B _13608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10750_ _10750_/A _10750_/B vssd1 vssd1 vccd1 vccd1 _10750_/X sky130_fd_sc_hd__or2_1
XFILLER_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10481__A1 _11099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09409_ _09409_/A vssd1 vssd1 vccd1 vccd1 _10219_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10681_ _09209_/A _10673_/X _10675_/X _10680_/X _10823_/A vssd1 vssd1 vccd1 vccd1
+ _10681_/X sky130_fd_sc_hd__a221o_1
X_12420_ _13712_/A vssd1 vssd1 vccd1 vccd1 _13702_/A sky130_fd_sc_hd__buf_2
XFILLER_138_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10769__C1 _09353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15848__S _15852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12351_ _09688_/A _18517_/Q _12423_/S vssd1 vssd1 vccd1 vccd1 _12372_/A sky130_fd_sc_hd__mux2_8
XFILLER_126_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10784__A2 _12469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11302_ _18421_/Q vssd1 vssd1 vccd1 vccd1 _14900_/A sky130_fd_sc_hd__clkbuf_2
X_15070_ _18489_/Q _15069_/B _14893_/A vssd1 vssd1 vccd1 vccd1 _15070_/X sky130_fd_sc_hd__a21o_1
X_12282_ _12282_/A vssd1 vssd1 vccd1 vccd1 _14253_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_153_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14021_ _11374_/A _11664_/A _11550_/B vssd1 vssd1 vccd1 vccd1 _14126_/A sky130_fd_sc_hd__a21o_4
XFILLER_107_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11233_ _11233_/A _11233_/B vssd1 vssd1 vccd1 vccd1 _11233_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09147__A _09147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10092__S0 _10153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11164_ _09689_/X _11155_/X _11159_/X _11163_/X _09134_/A vssd1 vssd1 vccd1 vccd1
+ _11164_/X sky130_fd_sc_hd__a311o_4
XFILLER_45_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10115_ _10115_/A _10115_/B vssd1 vssd1 vccd1 vccd1 _10115_/X sky130_fd_sc_hd__and2_1
XFILLER_1_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18760_ _19442_/CLK _18760_/D vssd1 vssd1 vccd1 vccd1 _18760_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13486__A1 _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15972_ _14761_/X _18986_/Q _15972_/S vssd1 vssd1 vccd1 vccd1 _15973_/A sky130_fd_sc_hd__mux2_1
X_11095_ _09434_/X _11086_/X _11090_/X _11094_/X _10373_/A vssd1 vssd1 vccd1 vccd1
+ _11095_/X sky130_fd_sc_hd__a311o_4
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_54_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19395_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17711_ _17711_/A vssd1 vssd1 vccd1 vccd1 _17711_/X sky130_fd_sc_hd__clkbuf_2
X_10046_ _19618_/Q _19456_/Q _18902_/Q _18672_/Q _09865_/A _10029_/A vssd1 vssd1 vccd1
+ vccd1 _10047_/B sky130_fd_sc_hd__mux4_1
XFILLER_29_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14923_ _14921_/X _14922_/X _14923_/S vssd1 vssd1 vccd1 vccd1 _14923_/X sky130_fd_sc_hd__mux2_1
X_18691_ _19633_/CLK _18691_/D vssd1 vssd1 vccd1 vccd1 _18691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output133_A _12462_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17642_ _13088_/A _17641_/Y _17658_/S vssd1 vssd1 vccd1 vccd1 _17642_/X sky130_fd_sc_hd__mux2_1
X_14854_ _11542_/X _14852_/X _14853_/X vssd1 vssd1 vccd1 vccd1 _16680_/A sky130_fd_sc_hd__o21a_4
XFILLER_36_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13805_ _13797_/X _13799_/Y _13800_/X _13804_/Y vssd1 vssd1 vccd1 vccd1 _13805_/X
+ sky130_fd_sc_hd__a31o_1
X_17573_ _19645_/Q _16797_/A _17579_/S vssd1 vssd1 vccd1 vccd1 _17574_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_69_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19818_/CLK sky130_fd_sc_hd__clkbuf_16
X_11997_ _11997_/A vssd1 vssd1 vccd1 vccd1 _11997_/X sky130_fd_sc_hd__buf_2
X_14785_ _14786_/A _14786_/C _18465_/Q vssd1 vssd1 vccd1 vccd1 _14787_/A sky130_fd_sc_hd__a21oi_1
X_19312_ _19539_/CLK _19312_/D vssd1 vssd1 vccd1 vccd1 _19312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16524_ _16524_/A vssd1 vssd1 vccd1 vccd1 _19219_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10948_ _10950_/A _10947_/X _10774_/X vssd1 vssd1 vccd1 vccd1 _10948_/X sky130_fd_sc_hd__o21a_1
X_13736_ _14120_/A vssd1 vssd1 vccd1 vccd1 _13736_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14738__A1 _14732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19243_ _19630_/CLK _19243_/D vssd1 vssd1 vccd1 vccd1 _19243_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10472__A1 _11099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16455_ _16501_/S vssd1 vssd1 vccd1 vccd1 _16464_/S sky130_fd_sc_hd__buf_4
XANTENNA__14738__B2 _14703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13667_ _13667_/A vssd1 vssd1 vccd1 vccd1 _13667_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10879_ _10864_/X _10869_/X _10878_/X _10823_/A vssd1 vssd1 vccd1 vccd1 _10879_/X
+ sky130_fd_sc_hd__a22o_1
X_15406_ _18750_/Q _15232_/X _15406_/S vssd1 vssd1 vccd1 vccd1 _15407_/A sky130_fd_sc_hd__mux2_1
X_12618_ _18338_/Q _12574_/X _12575_/X _12617_/X vssd1 vssd1 vccd1 vccd1 _18338_/D
+ sky130_fd_sc_hd__a31o_1
X_19174_ _19643_/CLK _19174_/D vssd1 vssd1 vccd1 vccd1 _19174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16386_ _16386_/A vssd1 vssd1 vccd1 vccd1 _19158_/D sky130_fd_sc_hd__clkbuf_1
X_13598_ _13598_/A vssd1 vssd1 vccd1 vccd1 _14192_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__17688__A0 _19674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18125_ _19828_/Q _18120_/C _18124_/Y vssd1 vssd1 vccd1 vccd1 _19828_/D sky130_fd_sc_hd__o21a_1
X_12549_ _12751_/B _12747_/C _12751_/D vssd1 vssd1 vccd1 vccd1 _12628_/A sky130_fd_sc_hd__or3_4
X_15337_ _18720_/Q _15238_/X _15337_/S vssd1 vssd1 vccd1 vccd1 _15338_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18056_ _19804_/Q _18053_/B _18055_/Y vssd1 vssd1 vccd1 vccd1 _19804_/D sky130_fd_sc_hd__o21a_1
XANTENNA__15163__A1 _15162_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15268_ _15324_/A vssd1 vssd1 vccd1 vccd1 _15337_/S sky130_fd_sc_hd__buf_6
XANTENNA__13174__B1 _13154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17007_ _17007_/A vssd1 vssd1 vccd1 vccd1 _19408_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15059__A _18488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14219_ _14150_/X _14056_/X _14218_/X _13823_/X vssd1 vssd1 vccd1 vccd1 _14219_/X
+ sky130_fd_sc_hd__a211o_1
X_15199_ _15199_/A vssd1 vssd1 vccd1 vccd1 _18669_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09760_ _10075_/S vssd1 vssd1 vccd1 vccd1 _09760_/X sky130_fd_sc_hd__clkbuf_4
X_18958_ _19414_/CLK _18958_/D vssd1 vssd1 vccd1 vccd1 _18958_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17909_ _17909_/A _17909_/B vssd1 vssd1 vccd1 vccd1 _17910_/A sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_115_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09691_ _10417_/S vssd1 vssd1 vccd1 vccd1 _09692_/A sky130_fd_sc_hd__clkbuf_4
X_18889_ _19444_/CLK _18889_/D vssd1 vssd1 vccd1 vccd1 _18889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_1_0_clock_A clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09528__S0 _10450_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12437__C1 _17711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10999__C1 _19695_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13042__A _13042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12204__A2 _14203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09125_ _09125_/A _18567_/Q vssd1 vssd1 vccd1 vccd1 _11339_/C sky130_fd_sc_hd__or2b_1
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13977__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11497__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10605__S _10605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16499__S _16501_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09958_ _09953_/Y _09956_/X _09957_/X _10042_/A vssd1 vssd1 vccd1 vccd1 _09958_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_131_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14958__D _14958_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _19526_/Q _19140_/Q _19590_/Q _18746_/Q _09803_/X _09810_/X vssd1 vssd1 vccd1
+ vccd1 _09890_/B sky130_fd_sc_hd__mux4_1
XANTENNA__14320__B _14324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ _11920_/A vssd1 vssd1 vccd1 vccd1 _11925_/A sky130_fd_sc_hd__clkinv_2
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _11851_/A _11901_/C vssd1 vssd1 vccd1 vccd1 _11851_/Y sky130_fd_sc_hd__nor2_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15090__A0 _18622_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12979__B1 _12922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _19633_/Q _19050_/Q _19087_/Q _18693_/Q _10719_/X _10772_/X vssd1 vssd1 vccd1
+ vccd1 _10803_/B sky130_fd_sc_hd__mux4_2
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _14570_/A _14572_/B vssd1 vssd1 vccd1 vccd1 _14570_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11782_ _11811_/A _13630_/A vssd1 vssd1 vccd1 vccd1 _11783_/B sky130_fd_sc_hd__nor2_1
XFILLER_13_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17906__A1 _12361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09430__A _09430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ _18592_/Q _19281_/Q _10733_/S vssd1 vssd1 vccd1 vccd1 _10733_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13521_ _13521_/A _13521_/B _13521_/C vssd1 vssd1 vccd1 vccd1 _13521_/X sky130_fd_sc_hd__and3_1
XFILLER_159_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16962__S _16964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13452_ _13452_/A vssd1 vssd1 vccd1 vccd1 _18386_/D sky130_fd_sc_hd__clkbuf_1
X_16240_ _16071_/X _19094_/Q _16246_/S vssd1 vssd1 vccd1 vccd1 _16241_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10664_ _18593_/Q _19282_/Q _10664_/S vssd1 vssd1 vccd1 vccd1 _10664_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12403_ _12403_/A _14308_/B vssd1 vssd1 vccd1 vccd1 _12404_/B sky130_fd_sc_hd__and2_1
XANTENNA__15578__S _15584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13383_ _18262_/Q _12582_/A _12584_/A _19851_/Q vssd1 vssd1 vccd1 vccd1 _13383_/X
+ sky130_fd_sc_hd__a22o_1
X_16171_ _16171_/A vssd1 vssd1 vccd1 vccd1 _19059_/D sky130_fd_sc_hd__clkbuf_1
X_10595_ _18826_/Q _19380_/Q _19542_/Q _18794_/Q _10579_/S _09514_/A vssd1 vssd1 vccd1
+ vccd1 _10596_/B sky130_fd_sc_hd__mux4_1
XFILLER_127_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10301__S1 _09555_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12334_ _19753_/Q _12335_/C _19754_/Q vssd1 vssd1 vccd1 vccd1 _12336_/A sky130_fd_sc_hd__a21oi_1
X_15122_ _18642_/Q _15116_/X _15118_/X _09951_/A vssd1 vssd1 vccd1 vccd1 _18642_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15053_ _14999_/X _15047_/X _15050_/Y _15052_/X vssd1 vssd1 vccd1 vccd1 _16734_/A
+ sky130_fd_sc_hd__a22o_4
X_12265_ _12265_/A _12265_/B vssd1 vssd1 vccd1 vccd1 _12265_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_147_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14004_ _14178_/A vssd1 vssd1 vccd1 vccd1 _14297_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11200__A _11200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11216_ _11472_/A _11282_/A _11285_/B vssd1 vssd1 vccd1 vccd1 _11216_/X sky130_fd_sc_hd__and3_1
X_19861_ _19861_/CLK _19861_/D vssd1 vssd1 vccd1 vccd1 _19861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12196_ _17628_/S vssd1 vssd1 vccd1 vccd1 _12196_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput82 _12142_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[18] sky130_fd_sc_hd__buf_2
X_18812_ _19643_/CLK _18812_/D vssd1 vssd1 vccd1 vccd1 _18812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11147_ _11147_/A vssd1 vssd1 vccd1 vccd1 _11149_/A sky130_fd_sc_hd__inv_2
Xoutput93 _12385_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[28] sky130_fd_sc_hd__buf_2
XFILLER_96_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19792_ _19795_/CLK _19792_/D vssd1 vssd1 vccd1 vccd1 _19792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18743_ _19838_/CLK _18743_/D vssd1 vssd1 vccd1 vccd1 _18743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15955_ _15955_/A vssd1 vssd1 vccd1 vccd1 _18978_/D sky130_fd_sc_hd__clkbuf_1
X_11078_ _11080_/B _11078_/B vssd1 vssd1 vccd1 vccd1 _11248_/C sky130_fd_sc_hd__nand2_1
X_10029_ _10029_/A vssd1 vssd1 vccd1 vccd1 _10029_/X sky130_fd_sc_hd__buf_2
XFILLER_64_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14906_ _14896_/X _14899_/Y _14905_/Y vssd1 vssd1 vccd1 vccd1 _16693_/A sky130_fd_sc_hd__a21oi_2
X_18674_ _19720_/CLK _18674_/D vssd1 vssd1 vccd1 vccd1 _18674_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12031__A _12057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10142__B1 _09414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15886_ _15886_/A vssd1 vssd1 vccd1 vccd1 _18946_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17625_ _19663_/Q _17624_/X _17625_/S vssd1 vssd1 vccd1 vccd1 _17626_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14959__A1 _18447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14837_ input3/X _14801_/X _14804_/X vssd1 vssd1 vccd1 vccd1 _14845_/A sky130_fd_sc_hd__a21oi_4
XFILLER_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12966__A _14673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15342__A _15410_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17556_ _17556_/A vssd1 vssd1 vccd1 vccd1 _19637_/D sky130_fd_sc_hd__clkbuf_1
X_14768_ _18431_/Q _13196_/B _14992_/S vssd1 vssd1 vccd1 vccd1 _14768_/X sky130_fd_sc_hd__mux2_2
XANTENNA__13631__A1 _12355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09340__A _10387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16507_ _16507_/A vssd1 vssd1 vccd1 vccd1 _19211_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10445__A1 _10219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13719_ _14285_/A _12510_/B _13927_/A vssd1 vssd1 vccd1 vccd1 _13719_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16872__S _16880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17487_ _17533_/S vssd1 vssd1 vccd1 vccd1 _17496_/S sky130_fd_sc_hd__buf_4
XFILLER_31_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14699_ _14699_/A vssd1 vssd1 vccd1 vccd1 _18585_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19226_ _19580_/CLK _19226_/D vssd1 vssd1 vccd1 vccd1 _19226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16438_ _16042_/X _19181_/Q _16442_/S vssd1 vssd1 vccd1 vccd1 _16439_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19157_ _19706_/CLK _19157_/D vssd1 vssd1 vccd1 vccd1 _19157_/Q sky130_fd_sc_hd__dfxtp_1
X_16369_ _19151_/Q _15503_/X _16369_/S vssd1 vssd1 vccd1 vccd1 _16370_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_41_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11945__A1 _12478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18108_ _17925_/B _18105_/B _18107_/Y vssd1 vssd1 vccd1 vccd1 _19823_/D sky130_fd_sc_hd__o21a_1
XFILLER_145_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19088_ _19635_/CLK _19088_/D vssd1 vssd1 vccd1 vccd1 _19088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18039_ _18170_/A vssd1 vssd1 vccd1 vccd1 _18039_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12370__A1 _12361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09812_ _09814_/A _09811_/X _09415_/X vssd1 vssd1 vccd1 vccd1 _09812_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10381__B1 _09708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09743_ _10127_/A _09743_/B vssd1 vssd1 vccd1 vccd1 _09743_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09674_ _09674_/A vssd1 vssd1 vccd1 vccd1 _09674_/Y sky130_fd_sc_hd__inv_2
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13471__S _13475_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11633__B1 _11940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10436__B2 _18438_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16782__S _16791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15398__S _15406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12728__A3 _12727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16083__A _16793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09108_ _11585_/B _11495_/B vssd1 vssd1 vccd1 vccd1 _09113_/A sky130_fd_sc_hd__or2_2
XANTENNA__15127__B2 _11222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10380_ _19611_/Q _19449_/Q _18895_/Q _18665_/Q _10417_/S _09554_/A vssd1 vssd1 vccd1
+ vccd1 _10380_/X sky130_fd_sc_hd__mux4_2
XFILLER_164_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13689__A1 _14111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12050_ _13295_/A _12075_/C vssd1 vssd1 vccd1 vccd1 _12050_/X sky130_fd_sc_hd__or2_1
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11001_ _10857_/X _10990_/X _10999_/X _11000_/Y vssd1 vssd1 vccd1 vccd1 _11619_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_89_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15861__S _15863_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12489__C _12489_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15740_ _15740_/A vssd1 vssd1 vccd1 vccd1 _18881_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12952_ _18294_/Q _18293_/Q _12952_/C vssd1 vssd1 vccd1 vccd1 _12957_/C sky130_fd_sc_hd__and3_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ _11899_/Y _11902_/Y _12016_/S vssd1 vssd1 vccd1 vccd1 _11903_/X sky130_fd_sc_hd__mux2_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _18851_/Q _15497_/X _15675_/S vssd1 vssd1 vccd1 vccd1 _15672_/A sky130_fd_sc_hd__mux2_1
X_12883_ _18274_/Q _12883_/B _12883_/C vssd1 vssd1 vccd1 vccd1 _12884_/C sky130_fd_sc_hd__and3_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _17410_/A vssd1 vssd1 vccd1 vccd1 _19572_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15162__A _16664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14622_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18390_ _19791_/CLK _18390_/D vssd1 vssd1 vccd1 vccd1 _18390_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _09927_/A _10799_/X _10809_/X _09306_/A _10810_/X vssd1 vssd1 vccd1 vccd1
+ _11834_/X sky130_fd_sc_hd__a32o_2
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17788__S _17794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17341_ _16774_/X _19542_/Q _17341_/S vssd1 vssd1 vccd1 vccd1 _17342_/A sky130_fd_sc_hd__mux2_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _18354_/Q _15255_/A vssd1 vssd1 vccd1 vccd1 _11767_/A sky130_fd_sc_hd__and2_1
X_14553_ _14553_/A _14559_/B vssd1 vssd1 vccd1 vccd1 _14553_/X sky130_fd_sc_hd__or2_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _18410_/Q _13387_/X _13508_/S vssd1 vssd1 vccd1 vccd1 _13505_/A sky130_fd_sc_hd__mux2_1
X_10716_ _10707_/Y _10714_/X _10715_/X _10701_/A vssd1 vssd1 vccd1 vccd1 _10716_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_17272_ _19511_/Q _16673_/X _17280_/S vssd1 vssd1 vccd1 vccd1 _17273_/A sky130_fd_sc_hd__mux2_1
X_11696_ _11696_/A vssd1 vssd1 vccd1 vccd1 _11696_/Y sky130_fd_sc_hd__inv_2
X_14484_ _14484_/A vssd1 vssd1 vccd1 vccd1 _18512_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19011_ _19592_/CLK _19011_/D vssd1 vssd1 vccd1 vccd1 _19011_/Q sky130_fd_sc_hd__dfxtp_1
X_16223_ _16223_/A vssd1 vssd1 vccd1 vccd1 _19086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13435_ _18650_/Q _13435_/B vssd1 vssd1 vccd1 vccd1 _13435_/X sky130_fd_sc_hd__or2_1
X_10647_ _11050_/S vssd1 vssd1 vccd1 vccd1 _10648_/S sky130_fd_sc_hd__buf_4
XFILLER_155_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13366_ _18375_/Q _13413_/B vssd1 vssd1 vccd1 vccd1 _13366_/X sky130_fd_sc_hd__or2_1
XFILLER_6_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16154_ _16154_/A vssd1 vssd1 vccd1 vccd1 _19051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11849__B _19735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10578_ _09274_/A _10568_/X _10577_/X _09281_/A _18435_/Q vssd1 vssd1 vccd1 vccd1
+ _10601_/B sky130_fd_sc_hd__a32o_4
XFILLER_115_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15105_ _18629_/Q _15102_/X _15104_/X _10554_/B vssd1 vssd1 vccd1 vccd1 _18629_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12317_ _19684_/Q _11989_/X _11790_/X vssd1 vssd1 vccd1 vccd1 _12317_/X sky130_fd_sc_hd__o21a_1
XFILLER_170_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13297_ _13297_/A vssd1 vssd1 vccd1 vccd1 _13297_/X sky130_fd_sc_hd__clkbuf_2
X_16085_ _16083_/X _19029_/Q _16097_/S vssd1 vssd1 vccd1 vccd1 _16086_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16721__A _16721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10038__S0 _09866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12248_ _19681_/Q _12390_/B vssd1 vssd1 vccd1 vccd1 _12248_/X sky130_fd_sc_hd__or2_1
X_15036_ input21/X _14960_/X _15000_/X vssd1 vssd1 vccd1 vccd1 _15036_/X sky130_fd_sc_hd__a21o_1
XFILLER_123_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17028__S _17036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19844_ _19851_/CLK _19844_/D vssd1 vssd1 vccd1 vccd1 _19844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12179_ _12181_/A _12180_/A vssd1 vssd1 vccd1 vccd1 _12182_/A sky130_fd_sc_hd__and2_1
XFILLER_96_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09335__A _18977_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19775_ _19858_/CLK _19775_/D vssd1 vssd1 vccd1 vccd1 _19775_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16867__S _16869_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16987_ _16987_/A vssd1 vssd1 vccd1 vccd1 _19400_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12104__B2 _12486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18726_ _19636_/CLK _18726_/D vssd1 vssd1 vccd1 vccd1 _18726_/Q sky130_fd_sc_hd__dfxtp_1
X_15938_ _15009_/X _18970_/Q _15946_/S vssd1 vssd1 vccd1 vccd1 _15939_/A sky130_fd_sc_hd__mux2_1
X_18657_ _19442_/CLK _18657_/D vssd1 vssd1 vccd1 vccd1 _18657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15869_ _15869_/A vssd1 vssd1 vccd1 vccd1 _18939_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10761__S1 _09482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17608_ _19467_/Q _14743_/A vssd1 vssd1 vccd1 vccd1 _17609_/B sky130_fd_sc_hd__or2b_1
XFILLER_92_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09390_ _09390_/A vssd1 vssd1 vccd1 vccd1 _09391_/A sky130_fd_sc_hd__buf_2
X_18588_ _19599_/CLK _18588_/D vssd1 vssd1 vccd1 vccd1 _18588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17539_ _17539_/A vssd1 vssd1 vccd1 vccd1 _19629_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11615__B1 _11614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09533__A1_N _18456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19209_ _19659_/CLK _19209_/D vssd1 vssd1 vccd1 vccd1 _19209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16107__S _16113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10944__A _10944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15011__S _15056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14317__C1 _14120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15946__S _15946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12343__A1 _19754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input1_A io_dbus_rdata[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09726_ _18875_/Q _19333_/Q _10125_/A vssd1 vssd1 vccd1 vccd1 _09727_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09657_ _09276_/A _09647_/X _09656_/X _09283_/A _18453_/Q vssd1 vssd1 vccd1 vccd1
+ _09688_/A sky130_fd_sc_hd__a32o_4
XFILLER_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _10451_/A vssd1 vssd1 vccd1 vccd1 _09735_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11550_ _14545_/A _11550_/B vssd1 vssd1 vccd1 vccd1 _11552_/B sky130_fd_sc_hd__nor2_1
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10501_ _10651_/A vssd1 vssd1 vccd1 vccd1 _10501_/X sky130_fd_sc_hd__buf_2
XFILLER_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11481_ _11360_/C _11481_/B vssd1 vssd1 vccd1 vccd1 _13520_/B sky130_fd_sc_hd__and2b_1
XFILLER_137_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13220_ _19768_/Q vssd1 vssd1 vccd1 vccd1 _17954_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10432_ _10432_/A _10432_/B vssd1 vssd1 vccd1 vccd1 _10432_/X sky130_fd_sc_hd__or2_1
XFILLER_148_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14045__B _14045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13151_ _13139_/X _13149_/X _13150_/X _13102_/X vssd1 vssd1 vccd1 vccd1 _18351_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10363_ _10910_/A vssd1 vssd1 vccd1 vccd1 _10364_/A sky130_fd_sc_hd__buf_2
XFILLER_151_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12102_ _17711_/A _12097_/X _12098_/X _12101_/X _11801_/X vssd1 vssd1 vccd1 vccd1
+ _12102_/X sky130_fd_sc_hd__a311o_1
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13082_ _19476_/Q _12669_/A _13428_/B _18390_/Q _13081_/X vssd1 vssd1 vccd1 vccd1
+ _13082_/X sky130_fd_sc_hd__a221o_1
XANTENNA_input57_A io_ibus_inst[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ _10288_/A _10293_/X _09681_/X vssd1 vssd1 vccd1 vccd1 _10294_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12334__A1 _19753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13531__B1 _13542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12033_ _10412_/A _18504_/Q _12060_/A vssd1 vssd1 vccd1 vccd1 _13607_/A sky130_fd_sc_hd__mux2_2
X_16910_ _16910_/A vssd1 vssd1 vccd1 vccd1 _19366_/D sky130_fd_sc_hd__clkbuf_1
X_17890_ _17890_/A _17890_/B vssd1 vssd1 vccd1 vccd1 _17891_/A sky130_fd_sc_hd__and2_1
XFILLER_132_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09155__A _10466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16841_ _16841_/A vssd1 vssd1 vccd1 vccd1 _16841_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14996__A _16822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16687__S _16687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10991__S1 _10960_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19560_ _19643_/CLK _19560_/D vssd1 vssd1 vccd1 vccd1 _19560_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_9_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16772_ _16771_/X _19315_/Q _16775_/S vssd1 vssd1 vccd1 vccd1 _16773_/A sky130_fd_sc_hd__mux2_1
X_13984_ _13984_/A _13984_/B vssd1 vssd1 vccd1 vccd1 _13984_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18511_ _18519_/CLK _18511_/D vssd1 vssd1 vccd1 vccd1 _18511_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15723_ _15723_/A vssd1 vssd1 vccd1 vccd1 _18874_/D sky130_fd_sc_hd__clkbuf_1
X_12935_ _12943_/A _12935_/B _12939_/C vssd1 vssd1 vccd1 vccd1 _18288_/D sky130_fd_sc_hd__nor3_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19491_ _19786_/CLK _19491_/D vssd1 vssd1 vccd1 vccd1 _19491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18618__D input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ _18818_/CLK _18442_/D vssd1 vssd1 vccd1 vccd1 _18442_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _18844_/Q _15577_/X _15658_/S vssd1 vssd1 vccd1 vccd1 _15655_/A sky130_fd_sc_hd__mux2_1
X_12866_ _12875_/D vssd1 vssd1 vccd1 vccd1 _12873_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _14624_/A _14605_/B vssd1 vssd1 vccd1 vccd1 _14606_/A sky130_fd_sc_hd__and2_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18373_ _18381_/CLK _18373_/D vssd1 vssd1 vccd1 vccd1 _18373_/Q sky130_fd_sc_hd__dfxtp_1
X_11817_ _12017_/B vssd1 vssd1 vccd1 vccd1 _11959_/B sky130_fd_sc_hd__clkbuf_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16138__D _16212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _15585_/A vssd1 vssd1 vccd1 vccd1 _18814_/D sky130_fd_sc_hd__clkbuf_1
X_12797_ _19866_/Q _19865_/Q _19864_/Q _18231_/C vssd1 vssd1 vccd1 vccd1 _18234_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_159_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17311__S _17313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17324_ _16749_/X _19534_/Q _17330_/S vssd1 vssd1 vccd1 vccd1 _17325_/A sky130_fd_sc_hd__mux2_1
X_14536_ _16919_/C _14522_/X _14533_/X _14535_/X vssd1 vssd1 vccd1 vccd1 _18531_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _11751_/B vssd1 vssd1 vccd1 vccd1 _11748_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10281__C1 _11119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17255_ _17255_/A vssd1 vssd1 vccd1 vccd1 _19503_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10764__A _10764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14467_ _14591_/B vssd1 vssd1 vccd1 vccd1 _14476_/S sky130_fd_sc_hd__clkbuf_2
X_11679_ _11678_/B _11827_/B _13166_/A vssd1 vssd1 vccd1 vccd1 _11679_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13140__A _13171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16206_ _16206_/A vssd1 vssd1 vccd1 vccd1 _19075_/D sky130_fd_sc_hd__clkbuf_1
X_13418_ _11406_/D _19499_/Q _13418_/S vssd1 vssd1 vccd1 vccd1 _13418_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17186_ _17186_/A vssd1 vssd1 vccd1 vccd1 _19482_/D sky130_fd_sc_hd__clkbuf_1
X_14398_ _14426_/A vssd1 vssd1 vccd1 vccd1 _14410_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_128_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16137_ _16919_/A _16357_/B _16919_/C vssd1 vssd1 vccd1 vccd1 _16213_/B sky130_fd_sc_hd__and3_1
XFILLER_6_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13349_ _18373_/Q _13352_/B vssd1 vssd1 vccd1 vccd1 _13349_/X sky130_fd_sc_hd__or2_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15511__A1 _15510_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16068_ _16135_/S vssd1 vssd1 vccd1 vccd1 _16081_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_88_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11128__A2 _11117_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15019_ _14875_/X _15016_/X _15017_/Y _15018_/Y _14898_/X vssd1 vssd1 vccd1 vccd1
+ _15019_/X sky130_fd_sc_hd__a221o_1
XFILLER_97_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19827_ _19866_/CLK _19827_/D vssd1 vssd1 vccd1 vccd1 _19827_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10431__S0 _09632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17282__A _17304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19758_ _19759_/CLK _19758_/D vssd1 vssd1 vccd1 vccd1 _19758_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13286__C1 _13285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09511_ _10712_/A vssd1 vssd1 vccd1 vccd1 _09512_/A sky130_fd_sc_hd__clkbuf_4
X_18709_ _19716_/CLK _18709_/D vssd1 vssd1 vccd1 vccd1 _18709_/Q sky130_fd_sc_hd__dfxtp_1
X_19689_ _19689_/CLK _19689_/D vssd1 vssd1 vccd1 vccd1 _19689_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_65_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09442_ _09538_/A vssd1 vssd1 vccd1 vccd1 _09442_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16775__A0 _16774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _18979_/Q vssd1 vssd1 vccd1 vccd1 _10695_/A sky130_fd_sc_hd__inv_2
XFILLER_12_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10811__B2 _10810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14069__A1 _18436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_163_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09709_ _09712_/A _09705_/X _09707_/X _09708_/X vssd1 vssd1 vccd1 vccd1 _09709_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10981_ _11026_/A _10981_/B vssd1 vssd1 vccd1 vccd1 _10981_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12720_ _18302_/Q _12564_/A _13222_/S _19481_/Q vssd1 vssd1 vccd1 vccd1 _12720_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16766__A0 _16765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12651_ _12651_/A vssd1 vssd1 vccd1 vccd1 _12651_/X sky130_fd_sc_hd__buf_2
XFILLER_31_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11602_ _11374_/A _11664_/A _11485_/A vssd1 vssd1 vccd1 vccd1 _11602_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_169_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12582_ _12582_/A vssd1 vssd1 vccd1 vccd1 _12582_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15370_ _15370_/A vssd1 vssd1 vccd1 vccd1 _18733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12783__B _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14321_ _11602_/Y _14324_/A _13797_/X _14320_/X vssd1 vssd1 vccd1 vccd1 _14321_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10263__C1 _09708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17191__A0 _18441_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11533_ _14513_/A _11298_/B vssd1 vssd1 vccd1 vccd1 _11534_/A sky130_fd_sc_hd__or2b_1
XFILLER_168_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17040_ _17040_/A vssd1 vssd1 vccd1 vccd1 _19423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11464_ _12658_/A _15241_/B vssd1 vssd1 vccd1 vccd1 _13442_/C sky130_fd_sc_hd__nor2_2
XFILLER_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14252_ _14088_/X _14249_/X _14251_/X vssd1 vssd1 vccd1 vccd1 _14252_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_99_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13203_ _13203_/A vssd1 vssd1 vccd1 vccd1 _13203_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10415_ _19255_/Q _19026_/Q _18957_/Q _19351_/Q _11087_/S _09142_/A vssd1 vssd1 vccd1
+ vccd1 _10416_/B sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_88_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11395_ _18545_/Q _18544_/Q _18543_/Q _18542_/Q vssd1 vssd1 vccd1 vccd1 _11413_/A
+ sky130_fd_sc_hd__or4_4
X_14183_ _13788_/A _14105_/Y _14182_/Y _14054_/A vssd1 vssd1 vccd1 vccd1 _14183_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13134_ _18619_/Q _13134_/B vssd1 vssd1 vccd1 vccd1 _13134_/X sky130_fd_sc_hd__or2_1
X_10346_ _09430_/A _10335_/X _10344_/X _09625_/X _10345_/Y vssd1 vssd1 vccd1 vccd1
+ _12483_/A sky130_fd_sc_hd__o32a_4
X_18991_ _19444_/CLK _18991_/D vssd1 vssd1 vccd1 vccd1 _18991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17942_ _18085_/A vssd1 vssd1 vccd1 vccd1 _17980_/A sky130_fd_sc_hd__buf_2
XFILLER_152_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13065_ _13067_/B _13067_/C _13064_/Y vssd1 vssd1 vccd1 vccd1 _18331_/D sky130_fd_sc_hd__o21a_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10277_ _18865_/Q _19323_/Q _10277_/S vssd1 vssd1 vccd1 vccd1 _10278_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12016_ _12013_/X _12015_/X _12016_/S vssd1 vssd1 vccd1 vccd1 _12016_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17873_ _17873_/A vssd1 vssd1 vccd1 vccd1 _19737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13533__A2_N _14565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16824_ _16824_/A vssd1 vssd1 vccd1 vccd1 _19331_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19612_ _19612_/CLK _19612_/D vssd1 vssd1 vccd1 vccd1 _19612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19543_ _19543_/CLK _19543_/D vssd1 vssd1 vccd1 vccd1 _19543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16755_ _16755_/A vssd1 vssd1 vccd1 vccd1 _16755_/X sky130_fd_sc_hd__clkbuf_2
X_13967_ _13965_/X _13966_/X _14085_/S vssd1 vssd1 vccd1 vccd1 _13967_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13283__A2 _13279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15706_ _18867_/Q _15548_/X _15708_/S vssd1 vssd1 vccd1 vccd1 _15707_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12918_ _12925_/C _12919_/C _18284_/Q vssd1 vssd1 vccd1 vccd1 _12920_/B sky130_fd_sc_hd__a21oi_1
X_19474_ _19689_/CLK _19474_/D vssd1 vssd1 vccd1 vccd1 _19474_/Q sky130_fd_sc_hd__dfxtp_1
X_16686_ _16686_/A vssd1 vssd1 vccd1 vccd1 _16686_/X sky130_fd_sc_hd__clkbuf_2
X_13898_ _13750_/X _13897_/X _13816_/X vssd1 vssd1 vccd1 vccd1 _13898_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18425_ _18509_/CLK _18425_/D vssd1 vssd1 vccd1 vccd1 _18425_/Q sky130_fd_sc_hd__dfxtp_1
X_15637_ _15637_/A vssd1 vssd1 vccd1 vccd1 _18836_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _12850_/B _12850_/C _18265_/Q vssd1 vssd1 vccd1 vccd1 _12851_/B sky130_fd_sc_hd__a21oi_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14232__A1 _12244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17041__S _17047_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18356_ _18357_/CLK _18356_/D vssd1 vssd1 vccd1 vccd1 _18356_/Q sky130_fd_sc_hd__dfxtp_1
X_15568_ _18809_/Q _15567_/X _15568_/S vssd1 vssd1 vccd1 vccd1 _15569_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17307_ _19527_/Q _16725_/X _17313_/S vssd1 vssd1 vccd1 vccd1 _17308_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17182__A0 _19481_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14519_ _14519_/A _14519_/B vssd1 vssd1 vccd1 vccd1 _14519_/X sky130_fd_sc_hd__or2_1
X_18287_ _19759_/CLK _18287_/D vssd1 vssd1 vccd1 vccd1 _18287_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_159_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10494__A _10494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16880__S _16880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15499_ _15499_/A vssd1 vssd1 vccd1 vccd1 _18787_/D sky130_fd_sc_hd__clkbuf_1
X_17238_ _18455_/Q _13412_/X _17241_/S vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__mux2_1
XFILLER_174_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17169_ _17169_/A vssd1 vssd1 vccd1 vccd1 _19477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09991_ _19523_/Q _19137_/Q _19587_/Q _18743_/Q _09983_/X _09984_/X vssd1 vssd1 vccd1
+ vccd1 _09992_/B sky130_fd_sc_hd__mux4_1
XFILLER_143_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10404__S0 _10224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10955__S1 _10910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16120__S _16129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10669__A _10669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10493__C1 _09681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09425_ _18578_/Q _11665_/B vssd1 vssd1 vccd1 vccd1 _09425_/Y sky130_fd_sc_hd__nor2_2
XFILLER_53_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12884__A _12904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09356_ _09501_/A vssd1 vssd1 vccd1 vccd1 _11113_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09287_ _19078_/Q vssd1 vssd1 vccd1 vccd1 _09624_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_165_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13734__B1 _14120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10200_ _18603_/Q _19292_/Q _10200_/S vssd1 vssd1 vccd1 vccd1 _10200_/X sky130_fd_sc_hd__mux2_1
X_11180_ _11180_/A _11180_/B vssd1 vssd1 vccd1 vccd1 _11180_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10131_ _18605_/Q _19294_/Q _10131_/S vssd1 vssd1 vccd1 vccd1 _10132_/B sky130_fd_sc_hd__mux2_1
XFILLER_121_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10062_ _09892_/A _10057_/X _10059_/X _10061_/X _09404_/A vssd1 vssd1 vccd1 vccd1
+ _10062_/X sky130_fd_sc_hd__a221o_1
XFILLER_48_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17126__S _17130_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14870_ input6/X _14801_/X _14804_/X vssd1 vssd1 vccd1 vccd1 _14877_/A sky130_fd_sc_hd__a21oi_2
XFILLER_75_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12778__B _12778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13821_ _13821_/A _14328_/B vssd1 vssd1 vccd1 vccd1 _13821_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09433__A _11205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16540_ _16540_/A vssd1 vssd1 vccd1 vccd1 _19226_/D sky130_fd_sc_hd__clkbuf_1
X_13752_ _13913_/S _13743_/X _13751_/X vssd1 vssd1 vccd1 vccd1 _13752_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10964_ _10973_/A _10963_/X _10827_/A vssd1 vssd1 vccd1 vccd1 _10964_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10298__B _12485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12703_ _12703_/A vssd1 vssd1 vccd1 vccd1 _12737_/A sky130_fd_sc_hd__clkbuf_2
X_16471_ _16090_/X _19196_/Q _16475_/S vssd1 vssd1 vccd1 vccd1 _16472_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13683_ _13681_/X _13682_/X _13768_/S vssd1 vssd1 vccd1 vccd1 _13683_/X sky130_fd_sc_hd__mux2_1
X_10895_ _10895_/A _10895_/B vssd1 vssd1 vccd1 vccd1 _10895_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18210_ _18210_/A _18210_/B vssd1 vssd1 vccd1 vccd1 _19857_/D sky130_fd_sc_hd__nor2_1
X_15422_ _18755_/Q _15146_/X _15426_/S vssd1 vssd1 vccd1 vccd1 _15423_/A sky130_fd_sc_hd__mux2_1
X_12634_ _13092_/S _12634_/B vssd1 vssd1 vccd1 vccd1 _12634_/X sky130_fd_sc_hd__and2b_1
X_19190_ _19223_/CLK _19190_/D vssd1 vssd1 vccd1 vccd1 _19190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18141_ _18165_/A _18141_/B _18141_/C vssd1 vssd1 vccd1 vccd1 _19833_/D sky130_fd_sc_hd__nor3_1
XFILLER_129_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17164__A0 _18433_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15353_ _15410_/S vssd1 vssd1 vccd1 vccd1 _15362_/S sky130_fd_sc_hd__buf_2
X_12565_ _13108_/A _13108_/B vssd1 vssd1 vccd1 vccd1 _15242_/C sky130_fd_sc_hd__or2_1
XFILLER_102_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14304_ _13832_/A _13901_/B _14012_/X vssd1 vssd1 vccd1 vccd1 _14304_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11203__A _11203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18072_ _19810_/Q _18069_/B _18071_/Y vssd1 vssd1 vccd1 vccd1 _19810_/D sky130_fd_sc_hd__o21a_1
X_11516_ _11516_/A vssd1 vssd1 vccd1 vccd1 _13524_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__10882__S0 _10724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15284_ _15284_/A vssd1 vssd1 vccd1 vccd1 _18695_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12496_ _12496_/A vssd1 vssd1 vccd1 vccd1 _12496_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_144_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09929__C1 _09826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17023_ _19416_/Q _16683_/X _17025_/S vssd1 vssd1 vccd1 vccd1 _17024_/A sky130_fd_sc_hd__mux2_1
X_14235_ _18448_/Q _14232_/X _14306_/S vssd1 vssd1 vccd1 vccd1 _14236_/A sky130_fd_sc_hd__mux2_1
X_11447_ _18345_/Q _18336_/Q _11720_/A vssd1 vssd1 vccd1 vccd1 _11447_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16205__S _16205_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14166_ _14320_/A _14168_/B _14092_/A _14165_/X vssd1 vssd1 vccd1 vccd1 _14166_/X
+ sky130_fd_sc_hd__o211a_1
X_11378_ _11479_/A _11481_/B _13521_/B _11378_/D vssd1 vssd1 vccd1 vccd1 _11610_/A
+ sky130_fd_sc_hd__and4b_1
XANTENNA_output88_A _12265_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13117_ _13354_/A vssd1 vssd1 vccd1 vccd1 _13311_/A sky130_fd_sc_hd__clkbuf_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _10329_/A _10328_/X vssd1 vssd1 vccd1 vccd1 _10329_/X sky130_fd_sc_hd__or2b_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _14097_/A vssd1 vssd1 vccd1 vccd1 _14097_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18974_ _19725_/CLK _18974_/D vssd1 vssd1 vccd1 vccd1 _18974_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ _19760_/Q _17925_/B _18105_/B vssd1 vssd1 vccd1 vccd1 _17926_/C sky130_fd_sc_hd__and3_1
X_13048_ _13058_/D vssd1 vssd1 vccd1 vccd1 _13055_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17036__S _17036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17856_ _17856_/A vssd1 vssd1 vccd1 vccd1 _19728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_1_0_clock_A clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16807_ _16806_/X _19326_/Q _16807_/S vssd1 vssd1 vccd1 vccd1 _16808_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09343__A _11188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17787_ _17787_/A vssd1 vssd1 vccd1 vccd1 _19696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14999_ _14999_/A vssd1 vssd1 vccd1 vccd1 _14999_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19526_ _19622_/CLK _19526_/D vssd1 vssd1 vccd1 vccd1 _19526_/Q sky130_fd_sc_hd__dfxtp_1
X_16738_ _19305_/Q _16737_/X _16741_/S vssd1 vssd1 vccd1 vccd1 _16739_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19457_ _19587_/CLK _19457_/D vssd1 vssd1 vccd1 vccd1 _19457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16669_ _16669_/A vssd1 vssd1 vccd1 vccd1 _19283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09210_ _09210_/A vssd1 vssd1 vccd1 vccd1 _09434_/A sky130_fd_sc_hd__clkbuf_2
X_18408_ _19788_/CLK _18408_/D vssd1 vssd1 vccd1 vccd1 _18408_/Q sky130_fd_sc_hd__dfxtp_1
X_19388_ _19452_/CLK _19388_/D vssd1 vssd1 vccd1 vccd1 _19388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11114__S1 _09483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ _09141_/A vssd1 vssd1 vccd1 vccd1 _09142_/A sky130_fd_sc_hd__buf_2
X_18339_ _18401_/CLK _18339_/D vssd1 vssd1 vccd1 vccd1 _18339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_111_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16904__A _16904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11113__A _11113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10625__S0 _10353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09974_ _18608_/Q _19297_/Q _10075_/S vssd1 vssd1 vccd1 vccd1 _09974_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15255__A _15255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12598__B _12598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09253__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_36_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13247__A2 _13245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16785__S _16791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17394__A0 _16743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09408_ _09408_/A vssd1 vssd1 vccd1 vccd1 _09409_/A sky130_fd_sc_hd__buf_2
X_10680_ _09179_/A _10679_/X _09224_/A vssd1 vssd1 vccd1 vccd1 _10680_/X sky130_fd_sc_hd__o21a_1
XFILLER_139_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12758__A1 _12757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09339_ _10579_/S vssd1 vssd1 vccd1 vccd1 _10387_/S sky130_fd_sc_hd__buf_4
XFILLER_40_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12350_ _14289_/A _12350_/B vssd1 vssd1 vccd1 vccd1 _12353_/A sky130_fd_sc_hd__xor2_1
XFILLER_166_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11301_ _11564_/A _12024_/A vssd1 vssd1 vccd1 vccd1 _14431_/C sky130_fd_sc_hd__or2_4
XFILLER_4_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12281_ _11148_/A _18514_/Q _12444_/S vssd1 vssd1 vccd1 vccd1 _12282_/A sky130_fd_sc_hd__mux2_8
XANTENNA__16025__S _16027_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09387__B1 _09320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14020_ _14086_/S _13998_/Y _13706_/A vssd1 vssd1 vccd1 vccd1 _14020_/X sky130_fd_sc_hd__a21o_1
X_11232_ _11234_/A _11230_/C _11230_/A vssd1 vssd1 vccd1 vccd1 _11233_/B sky130_fd_sc_hd__a21oi_1
XFILLER_153_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09428__A _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11163_ _11166_/A _11160_/X _11162_/X _09708_/X vssd1 vssd1 vccd1 vccd1 _11163_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10114_ _18868_/Q _19326_/Q _10114_/S vssd1 vssd1 vccd1 vccd1 _10115_/B sky130_fd_sc_hd__mux2_1
XFILLER_110_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15971_ _15971_/A vssd1 vssd1 vccd1 vccd1 _18985_/D sky130_fd_sc_hd__clkbuf_1
X_11094_ _09463_/A _11091_/X _11093_/X _09227_/A vssd1 vssd1 vccd1 vccd1 _11094_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_150_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17710_ _18477_/Q _17710_/B vssd1 vssd1 vccd1 vccd1 _17710_/Y sky130_fd_sc_hd__nand2_1
X_10045_ _18838_/Q _19392_/Q _19554_/Q _18806_/Q _09866_/A _10029_/X vssd1 vssd1 vccd1
+ vccd1 _10045_/X sky130_fd_sc_hd__mux4_1
XANTENNA__15165__A _16667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14922_ _18444_/Q _12615_/B _14922_/S vssd1 vssd1 vccd1 vccd1 _14922_/X sky130_fd_sc_hd__mux2_1
X_18690_ _19630_/CLK _18690_/D vssd1 vssd1 vccd1 vccd1 _18690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09163__A _09163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17641_ _17649_/C _17641_/B vssd1 vssd1 vccd1 vccd1 _17641_/Y sky130_fd_sc_hd__nand2_2
X_14853_ input4/X _14801_/X _14804_/X vssd1 vssd1 vccd1 vccd1 _14853_/X sky130_fd_sc_hd__a21o_1
XFILLER_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14435__A1 _19728_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13804_ _13839_/S _13800_/B _14092_/A vssd1 vssd1 vccd1 vccd1 _13804_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_63_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17572_ _17572_/A vssd1 vssd1 vccd1 vccd1 _19644_/D sky130_fd_sc_hd__clkbuf_1
X_14784_ _14784_/A vssd1 vssd1 vccd1 vccd1 _18592_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11996_ _13265_/A _12020_/C _17730_/A vssd1 vssd1 vccd1 vccd1 _11996_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19311_ _19537_/CLK _19311_/D vssd1 vssd1 vccd1 vccd1 _19311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16523_ _19219_/Q _15516_/X _16525_/S vssd1 vssd1 vccd1 vccd1 _16524_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10457__C1 _09393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13735_ _11046_/A _13566_/X _13731_/X _13734_/X vssd1 vssd1 vccd1 vccd1 _18426_/D
+ sky130_fd_sc_hd__a22o_1
X_10947_ _19632_/Q _19049_/Q _19086_/Q _18692_/Q _10719_/X _10772_/X vssd1 vssd1 vccd1
+ vccd1 _10947_/X sky130_fd_sc_hd__mux4_2
XFILLER_91_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09862__A1 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13413__A _18379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19242_ _19806_/CLK _19242_/D vssd1 vssd1 vccd1 vccd1 _19242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16454_ _16454_/A vssd1 vssd1 vccd1 vccd1 _19188_/D sky130_fd_sc_hd__clkbuf_1
X_13666_ _12401_/A _13665_/X _13668_/S vssd1 vssd1 vccd1 vccd1 _13666_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14738__A2 _14736_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10878_ _09209_/A _10871_/Y _10873_/Y _10875_/Y _10877_/Y vssd1 vssd1 vccd1 vccd1
+ _10878_/X sky130_fd_sc_hd__o32a_1
X_15405_ _15405_/A vssd1 vssd1 vccd1 vccd1 _18749_/D sky130_fd_sc_hd__clkbuf_1
X_12617_ _13092_/S _12617_/B vssd1 vssd1 vccd1 vccd1 _12617_/X sky130_fd_sc_hd__and2b_1
X_19173_ _19625_/CLK _19173_/D vssd1 vssd1 vccd1 vccd1 _19173_/Q sky130_fd_sc_hd__dfxtp_1
X_16385_ _19158_/Q _15526_/X _16391_/S vssd1 vssd1 vccd1 vccd1 _16386_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13597_ _14111_/A _14176_/B _13682_/S vssd1 vssd1 vccd1 vccd1 _13597_/X sky130_fd_sc_hd__mux2_1
X_18124_ _18159_/A _18131_/C vssd1 vssd1 vccd1 vccd1 _18124_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15336_ _15336_/A vssd1 vssd1 vccd1 vccd1 _18719_/D sky130_fd_sc_hd__clkbuf_1
X_12548_ _18340_/Q _12531_/Y _12543_/X _12547_/X vssd1 vssd1 vccd1 vccd1 _12548_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_157_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18055_ _18071_/A _18059_/C vssd1 vssd1 vccd1 vccd1 _18055_/Y sky130_fd_sc_hd__nor2_1
X_15267_ _16847_/B _17535_/A vssd1 vssd1 vccd1 vccd1 _15324_/A sky130_fd_sc_hd__nor2_4
XFILLER_145_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12479_ _12479_/A vssd1 vssd1 vccd1 vccd1 _12479_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13174__A1 _19663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17006_ _19408_/Q _16657_/X _17014_/S vssd1 vssd1 vccd1 vccd1 _17007_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09338__A _10836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14218_ _13795_/X _14213_/X _14215_/Y _14217_/X vssd1 vssd1 vccd1 vccd1 _14218_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15198_ _18669_/Q _15197_/X _15201_/S vssd1 vssd1 vccd1 vccd1 _15199_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15774__S _15780_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14149_ _18441_/Q _14120_/X _14148_/X vssd1 vssd1 vccd1 vccd1 _18441_/D sky130_fd_sc_hd__o21a_1
XFILLER_140_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18957_ _19609_/CLK _18957_/D vssd1 vssd1 vccd1 vccd1 _18957_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12699__A _14648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14674__B2 _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17908_ _17908_/A vssd1 vssd1 vccd1 vccd1 _19756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09690_ _11171_/A vssd1 vssd1 vccd1 vccd1 _11168_/A sky130_fd_sc_hd__buf_2
X_18888_ _19442_/CLK _18888_/D vssd1 vssd1 vccd1 vccd1 _18888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17839_ _17839_/A vssd1 vssd1 vccd1 vccd1 _19720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10160__A1 _09996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15623__A0 _18830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09528__S1 _09587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09302__B1 _15412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19509_ _19571_/CLK _19509_/D vssd1 vssd1 vccd1 vccd1 _19509_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_4_5_0_clock_A clkbuf_4_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14138__B _14138_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09124_ _11343_/C vssd1 vssd1 vccd1 vccd1 _11484_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13469__S _13475_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11497__B _18565_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09248__A _09248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09464__S0 _10350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17465__A _17533_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09957_ _19265_/Q _19036_/Q _18967_/Q _19361_/Q _09866_/A _09869_/A vssd1 vssd1 vccd1
+ vccd1 _09957_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_183_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19639_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__14665__B2 input47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09888_ _09944_/A _09888_/B vssd1 vssd1 vccd1 vccd1 _09888_/Y sky130_fd_sc_hd__nor2_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _11850_/A vssd1 vssd1 vccd1 vccd1 _11901_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _10946_/A _10801_/B vssd1 vssd1 vccd1 vccd1 _10801_/X sky130_fd_sc_hd__or2_1
XFILLER_54_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11100__A0 _18830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _11811_/A _13630_/A vssd1 vssd1 vccd1 vccd1 _11783_/A sky130_fd_sc_hd__and2_1
XFILLER_54_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10857__A _10857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13520_ _13520_/A _13520_/B _13520_/C vssd1 vssd1 vccd1 vccd1 _13521_/C sky130_fd_sc_hd__and3_1
X_10732_ _10732_/A vssd1 vssd1 vccd1 vccd1 _12469_/A sky130_fd_sc_hd__inv_2
XFILLER_158_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_121_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19481_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15859__S _15863_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13451_ _18386_/Q _13112_/A _13453_/S vssd1 vssd1 vccd1 vccd1 _13452_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10663_ _10663_/A vssd1 vssd1 vccd1 vccd1 _10664_/S sky130_fd_sc_hd__buf_4
XFILLER_40_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12402_ _12403_/A _14308_/B vssd1 vssd1 vccd1 vccd1 _12428_/A sky130_fd_sc_hd__nor2_1
X_16170_ _16077_/X _19059_/Q _16172_/S vssd1 vssd1 vccd1 vccd1 _16171_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13382_ _19496_/Q _12741_/X _13380_/X _13381_/X vssd1 vssd1 vccd1 vccd1 _13382_/X
+ sky130_fd_sc_hd__a211o_1
X_10594_ _19606_/Q _19444_/Q _18890_/Q _18660_/Q _09522_/A _09515_/A vssd1 vssd1 vccd1
+ vccd1 _10594_/X sky130_fd_sc_hd__mux4_1
X_15121_ _18641_/Q _15116_/X _15118_/X _10003_/B vssd1 vssd1 vccd1 vccd1 _18641_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11688__A _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12333_ _12371_/B _12333_/B vssd1 vssd1 vccd1 vccd1 _12333_/X sky130_fd_sc_hd__xor2_4
XFILLER_154_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_136_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19695_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15052_ _14744_/X _15051_/X _14842_/A vssd1 vssd1 vccd1 vccd1 _15052_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09158__A _11157_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12264_ _12233_/A _14227_/B _12241_/A vssd1 vssd1 vccd1 vccd1 _12265_/B sky130_fd_sc_hd__o21a_1
XFILLER_5_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09455__S0 _10465_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14003_ _14003_/A vssd1 vssd1 vccd1 vccd1 _14003_/X sky130_fd_sc_hd__buf_2
XANTENNA__11200__B _12503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11215_ _11475_/A _11484_/A _11296_/C vssd1 vssd1 vccd1 vccd1 _11285_/B sky130_fd_sc_hd__and3_1
X_19860_ _19861_/CLK _19860_/D vssd1 vssd1 vccd1 vccd1 _19860_/Q sky130_fd_sc_hd__dfxtp_1
X_12195_ _12715_/B vssd1 vssd1 vccd1 vccd1 _17628_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_96_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18811_ _19559_/CLK _18811_/D vssd1 vssd1 vccd1 vccd1 _18811_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput83 _12163_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[19] sky130_fd_sc_hd__buf_2
X_11146_ _11269_/A _11269_/B _11269_/C _11272_/A _11145_/Y vssd1 vssd1 vccd1 vccd1
+ _11225_/C sky130_fd_sc_hd__a311o_1
X_19791_ _19791_/CLK _19791_/D vssd1 vssd1 vccd1 vccd1 _19791_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput94 _12407_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[29] sky130_fd_sc_hd__buf_2
XANTENNA__14511__B _14519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18742_ _19818_/CLK _18742_/D vssd1 vssd1 vccd1 vccd1 _18742_/Q sky130_fd_sc_hd__dfxtp_1
X_11077_ _11077_/A _12473_/A vssd1 vssd1 vccd1 vccd1 _11078_/B sky130_fd_sc_hd__or2_1
X_15954_ _17779_/A _15954_/B vssd1 vssd1 vccd1 vccd1 _15955_/A sky130_fd_sc_hd__and2_2
XFILLER_163_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10028_ _09278_/A _10018_/X _10027_/X _09285_/A _18447_/Q vssd1 vssd1 vccd1 vccd1
+ _10051_/A sky130_fd_sc_hd__a32o_4
XFILLER_76_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14905_ input8/X _14901_/X _14904_/X vssd1 vssd1 vccd1 vccd1 _14905_/Y sky130_fd_sc_hd__a21oi_1
X_18673_ _19587_/CLK _18673_/D vssd1 vssd1 vccd1 vccd1 _18673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15885_ _14729_/X _18946_/Q _15891_/S vssd1 vssd1 vccd1 vccd1 _15886_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17624_ _13182_/X _17623_/Y _17628_/S vssd1 vssd1 vccd1 vccd1 _17624_/X sky130_fd_sc_hd__mux2_1
X_14836_ _14836_/A vssd1 vssd1 vccd1 vccd1 _18596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09621__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13092__A0 _13110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11870__B _13617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17555_ _19637_/Q _16771_/A _17557_/S vssd1 vssd1 vccd1 vccd1 _17556_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14767_ _15060_/B vssd1 vssd1 vccd1 vccd1 _14992_/S sky130_fd_sc_hd__clkbuf_2
X_11979_ _11979_/A vssd1 vssd1 vccd1 vccd1 _11980_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16506_ _19211_/Q _15487_/X _16514_/S vssd1 vssd1 vccd1 vccd1 _16507_/A sky130_fd_sc_hd__mux2_1
X_13718_ _13974_/A vssd1 vssd1 vccd1 vccd1 _13927_/A sky130_fd_sc_hd__clkbuf_2
X_17486_ _17486_/A vssd1 vssd1 vccd1 vccd1 _19606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14698_ _17890_/A _14698_/B vssd1 vssd1 vccd1 vccd1 _14699_/A sky130_fd_sc_hd__and2_1
XANTENNA__15769__S _15769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19225_ _19640_/CLK _19225_/D vssd1 vssd1 vccd1 vccd1 _19225_/Q sky130_fd_sc_hd__dfxtp_1
X_16437_ _16437_/A vssd1 vssd1 vccd1 vccd1 _19180_/D sky130_fd_sc_hd__clkbuf_1
X_13649_ _13811_/A _13648_/X _13743_/S vssd1 vssd1 vccd1 vccd1 _13649_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19156_ _19726_/CLK _19156_/D vssd1 vssd1 vccd1 vccd1 _19156_/Q sky130_fd_sc_hd__dfxtp_1
X_16368_ _16368_/A vssd1 vssd1 vccd1 vccd1 _19150_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18107_ _17925_/B _18105_/B _18082_/X vssd1 vssd1 vccd1 vccd1 _18107_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_145_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15319_ _15319_/A vssd1 vssd1 vccd1 vccd1 _18711_/D sky130_fd_sc_hd__clkbuf_1
X_19087_ _19540_/CLK _19087_/D vssd1 vssd1 vccd1 vccd1 _19087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10706__S _10706_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16299_ _16051_/X _19120_/Q _16307_/S vssd1 vssd1 vccd1 vccd1 _16300_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13147__A1 _19761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18038_ _19798_/Q _18033_/B _18037_/Y vssd1 vssd1 vccd1 vccd1 _19798_/D sky130_fd_sc_hd__o21a_1
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11158__B1 _09184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09997__S1 _09984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10007__A _10007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09811_ _19653_/Q _19070_/Q _19107_/Q _18713_/Q _09809_/X _09810_/X vssd1 vssd1 vccd1
+ vccd1 _09811_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10381__A1 _09640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09742_ _19527_/Q _19141_/Q _19591_/Q _18747_/Q _09734_/X _10186_/A vssd1 vssd1 vccd1
+ vccd1 _09743_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12222__A _18371_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10133__A1 _10132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ _18876_/Q _19334_/Q _09673_/S vssd1 vssd1 vccd1 vccd1 _09674_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13083__B1 _12628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10436__A2 _10426_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10841__C1 _10774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19720_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10819__S0 _10905_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09107_ _09107_/A vssd1 vssd1 vccd1 vccd1 _11528_/A sky130_fd_sc_hd__buf_2
XFILLER_108_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17907__B _17907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_68_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19812_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14612__A _14612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11000_ _18427_/Q _11046_/B vssd1 vssd1 vccd1 vccd1 _11000_/Y sky130_fd_sc_hd__nand2_1
XFILLER_131_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13228__A _18627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _18293_/Q _12952_/C _18294_/Q vssd1 vssd1 vccd1 vccd1 _12953_/B sky130_fd_sc_hd__a21oi_1
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14758__S _14923_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10124__B2 _18445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _11902_/A _11984_/D vssd1 vssd1 vccd1 vccd1 _11902_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17134__S _17134_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15670_ _15670_/A vssd1 vssd1 vccd1 vccd1 _18850_/D sky130_fd_sc_hd__clkbuf_1
X_12882_ _12883_/B _12883_/C _18274_/Q vssd1 vssd1 vccd1 vccd1 _12884_/B sky130_fd_sc_hd__a21oi_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15063__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _14621_/A vssd1 vssd1 vccd1 vccd1 _18561_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11833_ _10732_/A _11831_/X _12023_/B _14580_/A vssd1 vssd1 vccd1 vccd1 _11939_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_73_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13074__B1 _13063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16973__S _16975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _17340_/A vssd1 vssd1 vccd1 vccd1 _19541_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _18537_/Q _14550_/X _14551_/Y _14548_/X vssd1 vssd1 vccd1 vccd1 _18537_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _11764_/A _11764_/B vssd1 vssd1 vccd1 vccd1 _15255_/A sky130_fd_sc_hd__nand2_2
XANTENNA__11003__A_N _09480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13503_ _13503_/A vssd1 vssd1 vccd1 vccd1 _18409_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _17317_/S vssd1 vssd1 vccd1 vccd1 _17280_/S sky130_fd_sc_hd__buf_4
XFILLER_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10715_ _19250_/Q _19021_/Q _18952_/Q _19346_/Q _10706_/S _09352_/A vssd1 vssd1 vccd1
+ vccd1 _10715_/X sky130_fd_sc_hd__mux4_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14483_ _18512_/Q _12246_/A _14487_/S vssd1 vssd1 vccd1 vccd1 _14484_/A sky130_fd_sc_hd__mux2_1
X_11695_ _11695_/A _13653_/A vssd1 vssd1 vccd1 vccd1 _11699_/A sky130_fd_sc_hd__xnor2_1
X_19010_ _19724_/CLK _19010_/D vssd1 vssd1 vccd1 vccd1 _19010_/Q sky130_fd_sc_hd__dfxtp_1
X_16222_ _16045_/X _19086_/Q _16224_/S vssd1 vssd1 vccd1 vccd1 _16223_/A sky130_fd_sc_hd__mux2_1
X_13434_ _17925_/B _12665_/X _12602_/X _18110_/B _13433_/X vssd1 vssd1 vccd1 vccd1
+ _13435_/B sky130_fd_sc_hd__a221o_4
XFILLER_174_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10646_ _11051_/S vssd1 vssd1 vccd1 vccd1 _11050_/S sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_5_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_158_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16153_ _16051_/X _19051_/Q _16161_/S vssd1 vssd1 vccd1 vccd1 _16154_/A sky130_fd_sc_hd__mux2_1
X_13365_ _13365_/A vssd1 vssd1 vccd1 vccd1 _13413_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__12307__A _12307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10577_ _10570_/X _10572_/X _10574_/X _10576_/X _09245_/A vssd1 vssd1 vccd1 vccd1
+ _10577_/X sky130_fd_sc_hd__a221o_2
XFILLER_127_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15104_ _15111_/A vssd1 vssd1 vccd1 vccd1 _15104_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12316_ _12313_/Y _12315_/Y _12452_/S vssd1 vssd1 vccd1 vccd1 _12316_/X sky130_fd_sc_hd__mux2_1
X_16084_ _16116_/A vssd1 vssd1 vccd1 vccd1 _16097_/S sky130_fd_sc_hd__buf_2
XFILLER_138_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13296_ _13267_/X _13294_/X _13295_/X _13282_/X vssd1 vssd1 vccd1 vccd1 _18364_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15035_ _15035_/A vssd1 vssd1 vccd1 vccd1 _18613_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17309__S _17313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10038__S1 _09869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12247_ _12119_/S _12245_/X _12246_/Y _11979_/A vssd1 vssd1 vccd1 vccd1 _12247_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_174_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19843_ _19851_/CLK _19843_/D vssd1 vssd1 vccd1 vccd1 _19843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12178_ _10098_/X _18510_/Q _12444_/S vssd1 vssd1 vccd1 vccd1 _12180_/A sky130_fd_sc_hd__mux2_8
XANTENNA__15826__A0 _14792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ _11130_/A _12481_/A vssd1 vssd1 vccd1 vccd1 _11131_/A sky130_fd_sc_hd__nor2_1
X_19774_ _19858_/CLK _19774_/D vssd1 vssd1 vccd1 vccd1 _19774_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16986_ _16838_/X _19400_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16987_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18725_ _19700_/CLK _18725_/D vssd1 vssd1 vccd1 vccd1 _18725_/Q sky130_fd_sc_hd__dfxtp_1
X_15937_ _15937_/A vssd1 vssd1 vccd1 vccd1 _15946_/S sky130_fd_sc_hd__buf_4
XFILLER_37_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15353__A _15410_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15868_ _15022_/X _18939_/Q _15874_/S vssd1 vssd1 vccd1 vccd1 _15869_/A sky130_fd_sc_hd__mux2_1
X_18656_ _19442_/CLK _18656_/D vssd1 vssd1 vccd1 vccd1 _18656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09351__A _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14819_ _14811_/X _14814_/X _14817_/Y _14818_/X vssd1 vssd1 vccd1 vccd1 _16670_/A
+ sky130_fd_sc_hd__o31a_2
X_17607_ _18460_/Q _19467_/Q vssd1 vssd1 vccd1 vccd1 _17621_/C sky130_fd_sc_hd__nand2b_2
XFILLER_64_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18587_ _19436_/CLK _18587_/D vssd1 vssd1 vccd1 vccd1 _18587_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16883__S _16891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15799_ _15799_/A vssd1 vssd1 vccd1 vccd1 _18908_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11615__A1 _12460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17538_ _19629_/Q _16743_/A _17546_/S vssd1 vssd1 vccd1 vccd1 _17539_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17469_ _17469_/A vssd1 vssd1 vccd1 vccd1 _19598_/D sky130_fd_sc_hd__clkbuf_1
X_19208_ _19725_/CLK _19208_/D vssd1 vssd1 vccd1 vccd1 _19208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19139_ _19427_/CLK _19139_/D vssd1 vssd1 vccd1 vccd1 _19139_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17503__A0 _19614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12217__A _19749_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11646__A_N _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16123__S _16129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15817__A0 _14753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14151__B _14155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09725_ _10177_/A _09725_/B vssd1 vssd1 vccd1 vccd1 _09725_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13482__S _13486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11791__A _19733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09656_ _09689_/A _09649_/X _09651_/X _09655_/X _09247_/A vssd1 vssd1 vccd1 vccd1
+ _09656_/X sky130_fd_sc_hd__a311o_4
XFILLER_55_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09587_ _09587_/A vssd1 vssd1 vccd1 vccd1 _10451_/A sky130_fd_sc_hd__buf_2
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12803__B1 _12802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10500_ _10500_/A vssd1 vssd1 vccd1 vccd1 _10500_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__10290__B1 _09412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11480_ _13526_/B _11474_/B _13520_/A _13521_/A vssd1 vssd1 vccd1 vccd1 _11538_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09658__S0 _09342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10431_ _18829_/Q _19383_/Q _19545_/Q _18797_/Q _09632_/A _10368_/X vssd1 vssd1 vccd1
+ vccd1 _10432_/B sky130_fd_sc_hd__mux4_1
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16822__A _16822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13150_ _18351_/Q _13183_/B vssd1 vssd1 vccd1 vccd1 _13150_/X sky130_fd_sc_hd__or2_1
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10362_ _10349_/X _10351_/X _10356_/X _10428_/A _09212_/A vssd1 vssd1 vccd1 vccd1
+ _10373_/B sky130_fd_sc_hd__o221a_1
XFILLER_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12101_ _13312_/A _12123_/C _12100_/Y vssd1 vssd1 vccd1 vccd1 _12101_/X sky130_fd_sc_hd__o21a_1
XFILLER_151_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13081_ _19666_/Q _12624_/A _13080_/X vssd1 vssd1 vccd1 vccd1 _13081_/X sky130_fd_sc_hd__a21o_1
XFILLER_3_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10293_ _19613_/Q _19451_/Q _18897_/Q _18667_/Q _09675_/S _11113_/A vssd1 vssd1 vccd1
+ vccd1 _10293_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09436__A _10905_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12032_ _14124_/A _12032_/B vssd1 vssd1 vccd1 vccd1 _12035_/A sky130_fd_sc_hd__xnor2_1
XFILLER_78_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15872__S _15874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16840_ _16840_/A vssd1 vssd1 vccd1 vccd1 _19336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16771_ _16771_/A vssd1 vssd1 vccd1 vccd1 _16771_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13983_ _13975_/X _13976_/Y _13981_/X _13982_/X vssd1 vssd1 vccd1 vccd1 _13983_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_59_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15722_ _18874_/Q _15570_/X _15730_/S vssd1 vssd1 vccd1 vccd1 _15723_/A sky130_fd_sc_hd__mux2_1
X_18510_ _18510_/CLK _18510_/D vssd1 vssd1 vccd1 vccd1 _18510_/Q sky130_fd_sc_hd__dfxtp_1
X_12934_ _12934_/A vssd1 vssd1 vccd1 vccd1 _12939_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ _19496_/CLK _19490_/D vssd1 vssd1 vccd1 vccd1 _19490_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_84_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15036__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09171__A _09171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15653_ _15653_/A vssd1 vssd1 vccd1 vccd1 _18843_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17799__S _17805_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18441_ _19078_/CLK _18441_/D vssd1 vssd1 vccd1 vccd1 _18441_/Q sky130_fd_sc_hd__dfxtp_4
X_12865_ _18269_/Q _18268_/Q _18267_/Q _12865_/D vssd1 vssd1 vccd1 vccd1 _12875_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _14511_/A _13106_/B _14603_/X input56/X vssd1 vssd1 vccd1 vccd1 _14605_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _18395_/CLK _18372_/D vssd1 vssd1 vccd1 vccd1 _18372_/Q sky130_fd_sc_hd__dfxtp_2
X_11816_ _11813_/Y _11815_/X _12389_/S vssd1 vssd1 vccd1 vccd1 _11816_/X sky130_fd_sc_hd__mux2_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11058__C1 _10944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _18814_/Q _15583_/X _15584_/S vssd1 vssd1 vccd1 vccd1 _15585_/A sky130_fd_sc_hd__mux2_1
X_12796_ _19863_/Q _19862_/Q _19861_/Q _18222_/C vssd1 vssd1 vccd1 vccd1 _18231_/C
+ sky130_fd_sc_hd__and4_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _17323_/A vssd1 vssd1 vccd1 vccd1 _19533_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _14585_/A vssd1 vssd1 vccd1 vccd1 _14535_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11747_/A _11747_/B vssd1 vssd1 vccd1 vccd1 _11751_/B sky130_fd_sc_hd__xor2_4
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17254_ _19503_/Q _16648_/X _17258_/S vssd1 vssd1 vccd1 vccd1 _17255_/A sky130_fd_sc_hd__mux2_1
X_14466_ _14466_/A vssd1 vssd1 vccd1 vccd1 _18504_/D sky130_fd_sc_hd__clkbuf_1
X_11678_ _13166_/A _11678_/B _11827_/B vssd1 vssd1 vccd1 vccd1 _11678_/X sky130_fd_sc_hd__or3_1
XFILLER_128_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16205_ _16128_/X _19075_/Q _16205_/S vssd1 vssd1 vccd1 vccd1 _16206_/A sky130_fd_sc_hd__mux2_1
X_13417_ _19689_/Q _12703_/A _13428_/B _18413_/Q _13416_/X vssd1 vssd1 vccd1 vccd1
+ _13417_/X sky130_fd_sc_hd__a221o_1
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12022__A1 _12043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13140__B _18620_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17185_ _19482_/Q _17184_/X _17189_/S vssd1 vssd1 vccd1 vccd1 _17186_/A sky130_fd_sc_hd__mux2_1
X_10629_ _09210_/A _10622_/X _10624_/X _10628_/X _09245_/A vssd1 vssd1 vccd1 vccd1
+ _10629_/X sky130_fd_sc_hd__a311o_2
XANTENNA__10256__S _10256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14397_ _18478_/Q vssd1 vssd1 vccd1 vccd1 _17716_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16136_ _16136_/A vssd1 vssd1 vccd1 vccd1 _19045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13348_ _13267_/X _13346_/X _13347_/X _13317_/X vssd1 vssd1 vccd1 vccd1 _18372_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17039__S _17047_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16067_ _16777_/A vssd1 vssd1 vccd1 vccd1 _16067_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13279_ _13217_/X _13269_/Y _13278_/X _13229_/X _18632_/Q vssd1 vssd1 vccd1 vccd1
+ _13279_/X sky130_fd_sc_hd__a32o_4
XFILLER_64_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09346__A _10033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11128__A3 _11126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15018_ _15018_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _15018_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16878__S _16880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19826_ _19866_/CLK _19826_/D vssd1 vssd1 vccd1 vccd1 _19826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19757_ _19759_/CLK _19757_/D vssd1 vssd1 vccd1 vccd1 _19757_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_111_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16969_ _16813_/X _19392_/Q _16975_/S vssd1 vssd1 vccd1 vccd1 _16970_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10004__B _12493_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09510_ _09522_/A vssd1 vssd1 vccd1 vccd1 _10450_/S sky130_fd_sc_hd__buf_4
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18708_ _19616_/CLK _18708_/D vssd1 vssd1 vccd1 vccd1 _18708_/Q sky130_fd_sc_hd__dfxtp_1
X_19688_ _19689_/CLK _19688_/D vssd1 vssd1 vccd1 vccd1 _19688_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12500__A _12500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09441_ _10422_/A vssd1 vssd1 vccd1 vccd1 _09538_/A sky130_fd_sc_hd__buf_2
XFILLER_37_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18639_ _19628_/CLK _18639_/D vssd1 vssd1 vccd1 vccd1 _18639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09372_ _18784_/Q _19013_/Q _18944_/Q _19242_/Q _09369_/S _09370_/A vssd1 vssd1 vccd1
+ vccd1 _09372_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10272__B1 _09988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16642__A _16741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11772__B1 _19732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15258__A _15262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16788__S _16791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_106_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09708_ _09708_/A vssd1 vssd1 vccd1 vccd1 _09708_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__12410__A _19757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10980_ _19244_/Q _19015_/Q _18946_/Q _19340_/Q _10663_/A _10364_/A vssd1 vssd1 vccd1
+ vccd1 _10981_/B sky130_fd_sc_hd__mux4_1
XFILLER_28_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09639_ _18780_/Q _19009_/Q _18940_/Q _19238_/Q _09643_/S _09695_/A vssd1 vssd1 vccd1
+ vccd1 _09640_/B sky130_fd_sc_hd__mux4_1
XFILLER_55_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14777__A0 _18432_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12650_ _18255_/Q vssd1 vssd1 vccd1 vccd1 _12821_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11601_ _09113_/B _11474_/B _13572_/B _11281_/Y vssd1 vssd1 vccd1 vccd1 _13587_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_169_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ _12603_/A vssd1 vssd1 vccd1 vccd1 _12582_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12783__C _15134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14320_ _14320_/A _14324_/B vssd1 vssd1 vccd1 vccd1 _14320_/X sky130_fd_sc_hd__or2_1
XFILLER_156_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11532_ _14543_/A _11333_/X _11476_/B _11531_/X _11378_/D vssd1 vssd1 vccd1 vccd1
+ _11538_/C sky130_fd_sc_hd__o311a_1
XFILLER_129_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17191__A1 _13307_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14251_ _14126_/A _12280_/A _13975_/A _14250_/Y vssd1 vssd1 vccd1 vccd1 _14251_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_137_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11463_ _11716_/A _11463_/B _11463_/C vssd1 vssd1 vccd1 vccd1 _15241_/B sky130_fd_sc_hd__nand3_2
XANTENNA__10076__S _10076_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13202_ _13248_/A _18625_/Q vssd1 vssd1 vccd1 vccd1 _13202_/Y sky130_fd_sc_hd__nand2_1
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10414_ _10414_/A vssd1 vssd1 vccd1 vccd1 _11262_/A sky130_fd_sc_hd__inv_2
Xclkbuf_opt_4_0_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_4_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_171_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14182_ _14182_/A _14182_/B vssd1 vssd1 vccd1 vccd1 _14182_/Y sky130_fd_sc_hd__nand2_1
X_11394_ _18551_/Q _18550_/Q _18553_/Q _18552_/Q vssd1 vssd1 vccd1 vccd1 _11400_/A
+ sky130_fd_sc_hd__or4bb_4
XFILLER_109_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11763__B1 _11720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13133_ _19760_/Q _13123_/X _13129_/X _13132_/X vssd1 vssd1 vccd1 vccd1 _13134_/B
+ sky130_fd_sc_hd__a211o_4
XANTENNA__15168__A _16670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10345_ _18441_/Q vssd1 vssd1 vccd1 vccd1 _10345_/Y sky130_fd_sc_hd__inv_2
X_18990_ _19541_/CLK _18990_/D vssd1 vssd1 vccd1 vccd1 _18990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13504__A1 _13387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17941_ _17944_/B _17944_/C _17940_/Y vssd1 vssd1 vccd1 vccd1 _19765_/D sky130_fd_sc_hd__o21a_1
X_13064_ _13067_/B _13067_/C _13063_/X vssd1 vssd1 vccd1 vccd1 _13064_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_112_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10276_ _10288_/A _10276_/B vssd1 vssd1 vccd1 vccd1 _10276_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10318__A1 _19194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12015_ _12043_/A _12067_/D vssd1 vssd1 vccd1 vccd1 _12015_/X sky130_fd_sc_hd__xor2_1
X_17872_ _17874_/A _17872_/B vssd1 vssd1 vccd1 vccd1 _17873_/A sky130_fd_sc_hd__or2_1
XFILLER_39_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1_0_clock_A clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19611_ _19708_/CLK _19611_/D vssd1 vssd1 vccd1 vccd1 _19611_/Q sky130_fd_sc_hd__dfxtp_1
X_16823_ _16822_/X _19331_/Q _16823_/S vssd1 vssd1 vccd1 vccd1 _16824_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19542_ _19639_/CLK _19542_/D vssd1 vssd1 vccd1 vccd1 _19542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12320__A _18375_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13966_ _13840_/X _13844_/X _13966_/S vssd1 vssd1 vccd1 vccd1 _13966_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16754_ _16754_/A vssd1 vssd1 vccd1 vccd1 _19309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12917_ _12991_/A vssd1 vssd1 vccd1 vccd1 _12943_/A sky130_fd_sc_hd__clkbuf_2
X_15705_ _15705_/A vssd1 vssd1 vccd1 vccd1 _18866_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19473_ _19791_/CLK _19473_/D vssd1 vssd1 vccd1 vccd1 _19473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16685_ _16685_/A vssd1 vssd1 vccd1 vccd1 _19288_/D sky130_fd_sc_hd__clkbuf_1
X_13897_ _13881_/S _13649_/X _13813_/Y vssd1 vssd1 vccd1 vccd1 _13897_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14768__A0 _18431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18424_ _19467_/CLK _18424_/D vssd1 vssd1 vccd1 vccd1 _18424_/Q sky130_fd_sc_hd__dfxtp_1
X_12848_ _12850_/B _12850_/C _12847_/Y vssd1 vssd1 vccd1 vccd1 _18264_/D sky130_fd_sc_hd__o21a_1
X_15636_ _18836_/Q _15551_/X _15636_/S vssd1 vssd1 vccd1 vccd1 _15637_/A sky130_fd_sc_hd__mux2_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13440__A0 _13112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15567_ _16822_/A vssd1 vssd1 vccd1 vccd1 _15567_/X sky130_fd_sc_hd__clkbuf_2
X_18355_ _18357_/CLK _18355_/D vssd1 vssd1 vccd1 vccd1 _18355_/Q sky130_fd_sc_hd__dfxtp_2
X_12779_ _12556_/X _12767_/Y _12778_/X _12712_/X _18643_/Q vssd1 vssd1 vccd1 vccd1
+ _12779_/X sky130_fd_sc_hd__a32o_4
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17306_ _17306_/A vssd1 vssd1 vccd1 vccd1 _19526_/D sky130_fd_sc_hd__clkbuf_1
X_14518_ _14518_/A vssd1 vssd1 vccd1 vccd1 _18526_/D sky130_fd_sc_hd__clkbuf_1
X_18286_ _19759_/CLK _18286_/D vssd1 vssd1 vccd1 vccd1 _18286_/Q sky130_fd_sc_hd__dfxtp_1
X_15498_ _18787_/Q _15497_/X _15504_/S vssd1 vssd1 vccd1 vccd1 _15499_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17237_ _17237_/A vssd1 vssd1 vccd1 vccd1 _19497_/D sky130_fd_sc_hd__clkbuf_1
X_14449_ _14449_/A vssd1 vssd1 vccd1 vccd1 _18496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17168_ _19477_/Q _17167_/X _17172_/S vssd1 vssd1 vccd1 vccd1 _17169_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16119_ _16829_/A vssd1 vssd1 vccd1 vccd1 _16119_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09990_ _09217_/A _09981_/X _09986_/X _09989_/X _09854_/A vssd1 vssd1 vccd1 vccd1
+ _09990_/X sky130_fd_sc_hd__a221o_2
X_17099_ _17121_/A vssd1 vssd1 vccd1 vccd1 _17108_/S sky130_fd_sc_hd__buf_4
XFILLER_170_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17293__A _17304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10404__S1 _11111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15248__A1 _17730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09804__A _09810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19809_ _19810_/CLK _19809_/D vssd1 vssd1 vccd1 vccd1 _19809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13326__A _18288_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12230__A _14227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10168__S0 _10076_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09424_ _09415_/X _09417_/Y _09419_/Y _09421_/Y _09423_/Y vssd1 vssd1 vccd1 vccd1
+ _09424_/X sky130_fd_sc_hd__o32a_1
XANTENNA__14759__B1 _14758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09355_ _10384_/A vssd1 vssd1 vccd1 vccd1 _09501_/A sky130_fd_sc_hd__buf_2
XANTENNA__13431__B1 _12703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09286_ _09233_/X _09250_/X _09278_/X _09285_/X _18457_/Q vssd1 vssd1 vccd1 vccd1
+ _11205_/A sky130_fd_sc_hd__a32o_4
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10340__S0 _10129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13996__A _13996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_32_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13734__A1 _12511_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10130_ _10130_/A vssd1 vssd1 vccd1 vccd1 _10130_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10061_ _10044_/A _10060_/X _09318_/A vssd1 vssd1 vccd1 vccd1 _10061_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17407__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09714__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13236__A _13236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13820_ _13810_/X _13817_/X _13819_/X vssd1 vssd1 vccd1 vccd1 _14328_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__09433__B _12505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13751_ _13745_/X _13748_/X _13750_/X vssd1 vssd1 vccd1 vccd1 _13751_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__13670__A0 _12446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10963_ _19632_/Q _19049_/Q _19086_/Q _18692_/Q _10663_/A _10364_/A vssd1 vssd1 vccd1
+ vccd1 _10963_/X sky130_fd_sc_hd__mux4_2
XFILLER_90_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13670__S _13724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12702_ _19867_/Q vssd1 vssd1 vccd1 vccd1 _18239_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16470_ _16470_/A vssd1 vssd1 vccd1 vccd1 _19195_/D sky130_fd_sc_hd__clkbuf_1
X_13682_ _13615_/Y _14045_/B _13682_/S vssd1 vssd1 vccd1 vccd1 _13682_/X sky130_fd_sc_hd__mux2_1
X_10894_ _19503_/Q _19117_/Q _19567_/Q _18723_/Q _10711_/A _10785_/X vssd1 vssd1 vccd1
+ vccd1 _10895_/B sky130_fd_sc_hd__mux4_2
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15421_ _15421_/A vssd1 vssd1 vccd1 vccd1 _18754_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12225__A1 _19749_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12633_ _12600_/X _12619_/Y _12632_/X _12558_/X _18638_/Q vssd1 vssd1 vccd1 vccd1
+ _12634_/B sky130_fd_sc_hd__a32o_4
XFILLER_54_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18140_ _19833_/Q _18140_/B _18140_/C vssd1 vssd1 vccd1 vccd1 _18141_/C sky130_fd_sc_hd__and3_1
X_15352_ _15352_/A vssd1 vssd1 vccd1 vccd1 _18725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12564_ _12564_/A vssd1 vssd1 vccd1 vccd1 _13108_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17164__A1 _13088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14303_ _13971_/X _13892_/X _14302_/X vssd1 vssd1 vccd1 vccd1 _14303_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15597__S _15603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18071_ _18071_/A _18075_/C vssd1 vssd1 vccd1 vccd1 _18071_/Y sky130_fd_sc_hd__nor2_1
X_11515_ _18575_/Q vssd1 vssd1 vccd1 vccd1 _14566_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15283_ _18695_/Q _15159_/X _15289_/S vssd1 vssd1 vccd1 vccd1 _15284_/A sky130_fd_sc_hd__mux2_1
X_12495_ _12495_/A _12495_/B _12495_/C vssd1 vssd1 vccd1 vccd1 _12496_/A sky130_fd_sc_hd__and3_1
XANTENNA__10882__S1 _10726_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17022_ _17022_/A vssd1 vssd1 vccd1 vccd1 _19415_/D sky130_fd_sc_hd__clkbuf_1
X_14234_ _14384_/A vssd1 vssd1 vccd1 vccd1 _14306_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__14922__A0 _18444_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11446_ _18348_/Q _18342_/Q _18382_/Q _18349_/Q vssd1 vssd1 vccd1 vccd1 _11720_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_125_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14165_ _14285_/A _14168_/A vssd1 vssd1 vccd1 vccd1 _14165_/X sky130_fd_sc_hd__or2_1
X_11377_ _11333_/X _13583_/A _11639_/A _11531_/A vssd1 vssd1 vccd1 vccd1 _11378_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_153_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13116_ _14431_/A _15242_/C _13119_/C vssd1 vssd1 vccd1 vccd1 _13354_/A sky130_fd_sc_hd__or3b_2
XFILLER_98_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ _18864_/Q _19322_/Q _10328_/S vssd1 vssd1 vccd1 vccd1 _10328_/X sky130_fd_sc_hd__mux2_1
X_18973_ _19271_/CLK _18973_/D vssd1 vssd1 vccd1 vccd1 _18973_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14096_ _14150_/A _14087_/X _14095_/X _13950_/X vssd1 vssd1 vccd1 vccd1 _14096_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12034__B _13607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17317__S _17317_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13845__S _13845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17924_ _17925_/B _18105_/B _19760_/Q vssd1 vssd1 vccd1 vccd1 _17926_/B sky130_fd_sc_hd__a21oi_1
X_13047_ _18326_/Q _18325_/Q _18327_/Q _13047_/D vssd1 vssd1 vccd1 vccd1 _13058_/D
+ sky130_fd_sc_hd__and4_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10259_ _09146_/A _10256_/X _10258_/X vssd1 vssd1 vccd1 vccd1 _10259_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17855_ _17895_/A _19728_/Q _17855_/C vssd1 vssd1 vccd1 vccd1 _17856_/A sky130_fd_sc_hd__and3_1
XFILLER_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16806_ _16806_/A vssd1 vssd1 vccd1 vccd1 _16806_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12050__A _13295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17786_ _15133_/X _19696_/Q _17794_/S vssd1 vssd1 vccd1 vccd1 _17787_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14998_ _14998_/A vssd1 vssd1 vccd1 vccd1 _18610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19525_ _19720_/CLK _19525_/D vssd1 vssd1 vccd1 vccd1 _19525_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13661__A0 _14289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16737_ _16737_/A vssd1 vssd1 vccd1 vccd1 _16737_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13949_ _13949_/A _13949_/B vssd1 vssd1 vccd1 vccd1 _13949_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_3_5_0_clock_A clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17052__S _17058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19456_ _19618_/CLK _19456_/D vssd1 vssd1 vccd1 vccd1 _19456_/Q sky130_fd_sc_hd__dfxtp_1
X_16668_ _19283_/Q _16667_/X _16671_/S vssd1 vssd1 vccd1 vccd1 _16669_/A sky130_fd_sc_hd__mux2_1
X_18407_ _19788_/CLK _18407_/D vssd1 vssd1 vccd1 vccd1 _18407_/Q sky130_fd_sc_hd__dfxtp_1
X_15619_ _18828_/Q _15526_/X _15625_/S vssd1 vssd1 vccd1 vccd1 _15620_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16891__S _16891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19387_ _19549_/CLK _19387_/D vssd1 vssd1 vccd1 vccd1 _19387_/Q sky130_fd_sc_hd__dfxtp_1
X_16599_ _19255_/Q vssd1 vssd1 vccd1 vccd1 _16600_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_148_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09140_ _10422_/A vssd1 vssd1 vccd1 vccd1 _09141_/A sky130_fd_sc_hd__clkbuf_2
X_18338_ _18401_/CLK _18338_/D vssd1 vssd1 vccd1 vccd1 _18338_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12209__B _14216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18269_ _19472_/CLK _18269_/D vssd1 vssd1 vccd1 vccd1 _18269_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15300__S _15300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09396__A1 _09320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10625__S1 _10548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09973_ _09927_/X _09963_/X _09972_/X _09309_/X _18448_/Q vssd1 vssd1 vccd1 vccd1
+ _12493_/C sky130_fd_sc_hd__a32o_4
XFILLER_58_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09534__A _11202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15970__S _15972_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09407_ _09407_/A vssd1 vssd1 vccd1 vccd1 _09408_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12207__A1 _10051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09338_ _10836_/A vssd1 vssd1 vccd1 vccd1 _10579_/S sky130_fd_sc_hd__buf_2
XANTENNA__17146__A1 _18428_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10769__A1 _10650_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ _14551_/A _16138_/B _09265_/Y _09267_/X _09268_/Y vssd1 vssd1 vccd1 vccd1
+ _11368_/C sky130_fd_sc_hd__o2111a_1
XFILLER_138_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11300_ _11575_/B vssd1 vssd1 vccd1 vccd1 _12024_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12280_ _12280_/A _12280_/B vssd1 vssd1 vccd1 vccd1 _12284_/A sky130_fd_sc_hd__xnor2_1
XFILLER_154_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09387__A1 _09814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11231_ _11229_/Y _11139_/X _10197_/A _11233_/A vssd1 vssd1 vccd1 vccd1 _11231_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11194__A1 _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11162_ _11171_/A _11162_/B vssd1 vssd1 vccd1 vccd1 _11162_/X sky130_fd_sc_hd__or2_1
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10113_ _19262_/Q _19033_/Q _18964_/Q _19358_/Q _10094_/X _10103_/X vssd1 vssd1 vccd1
+ vccd1 _10113_/X sky130_fd_sc_hd__mux4_1
X_15970_ _14753_/X _18985_/Q _15972_/S vssd1 vssd1 vccd1 vccd1 _15971_/A sky130_fd_sc_hd__mux2_1
X_11093_ _11102_/A _11093_/B vssd1 vssd1 vccd1 vccd1 _11093_/X sky130_fd_sc_hd__or2_1
XFILLER_103_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12143__B1 _19746_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input32_A io_dbus_rdata[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09444__A _11097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ _10044_/A _10044_/B vssd1 vssd1 vccd1 vccd1 _10044_/X sky130_fd_sc_hd__or2_1
X_14921_ _17701_/B _14932_/C vssd1 vssd1 vccd1 vccd1 _14921_/X sky130_fd_sc_hd__xor2_1
XFILLER_102_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17082__A0 _16768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17640_ _18465_/Q _17640_/B vssd1 vssd1 vccd1 vccd1 _17641_/B sky130_fd_sc_hd__nand2_1
XFILLER_75_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14852_ _14850_/X _14851_/X _14945_/B vssd1 vssd1 vccd1 vccd1 _14852_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13803_ _14088_/A vssd1 vssd1 vccd1 vccd1 _14092_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14783_ _14782_/X _18592_/Q _14822_/S vssd1 vssd1 vccd1 vccd1 _14784_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17571_ _19644_/Q _16793_/A _17579_/S vssd1 vssd1 vccd1 vccd1 _17572_/A sky130_fd_sc_hd__mux2_1
X_11995_ _12091_/A vssd1 vssd1 vccd1 vccd1 _17730_/A sky130_fd_sc_hd__buf_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19310_ _19691_/CLK _19310_/D vssd1 vssd1 vccd1 vccd1 _19310_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15181__A _16683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16522_ _16522_/A vssd1 vssd1 vccd1 vccd1 _19218_/D sky130_fd_sc_hd__clkbuf_1
X_13734_ _12511_/Y _13933_/A _14120_/A vssd1 vssd1 vccd1 vccd1 _13734_/X sky130_fd_sc_hd__o21a_1
X_10946_ _10946_/A _10946_/B vssd1 vssd1 vccd1 vccd1 _10946_/X sky130_fd_sc_hd__or2_1
XFILLER_44_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19241_ _19337_/CLK _19241_/D vssd1 vssd1 vccd1 vccd1 _19241_/Q sky130_fd_sc_hd__dfxtp_1
X_13665_ _13665_/A vssd1 vssd1 vccd1 vccd1 _13665_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16453_ _16064_/X _19188_/Q _16453_/S vssd1 vssd1 vccd1 vccd1 _16454_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14738__A3 _14737_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10877_ _10871_/A _10876_/X _10827_/X vssd1 vssd1 vccd1 vccd1 _10877_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15404_ _18749_/Q _15229_/X _15406_/S vssd1 vssd1 vccd1 vccd1 _15405_/A sky130_fd_sc_hd__mux2_1
X_12616_ _12600_/X _12601_/Y _12615_/X _12558_/X _18637_/Q vssd1 vssd1 vccd1 vccd1
+ _12617_/B sky130_fd_sc_hd__a32o_4
X_19172_ _19721_/CLK _19172_/D vssd1 vssd1 vccd1 vccd1 _19172_/Q sky130_fd_sc_hd__dfxtp_1
X_16384_ _16384_/A vssd1 vssd1 vccd1 vccd1 _19157_/D sky130_fd_sc_hd__clkbuf_1
X_13596_ _13596_/A vssd1 vssd1 vccd1 vccd1 _14176_/B sky130_fd_sc_hd__buf_2
XANTENNA__10304__S0 _09553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18123_ _18133_/D vssd1 vssd1 vccd1 vccd1 _18131_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15335_ _18719_/Q _15235_/X _15337_/S vssd1 vssd1 vccd1 vccd1 _15336_/A sky130_fd_sc_hd__mux2_1
X_12547_ _18283_/Q _13156_/A _12642_/A _13312_/A vssd1 vssd1 vccd1 vccd1 _12547_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16216__S _16224_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18054_ _18054_/A vssd1 vssd1 vccd1 vccd1 _18059_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15266_ _16430_/A _16919_/B _15412_/C vssd1 vssd1 vccd1 vccd1 _17535_/A sky130_fd_sc_hd__or3b_4
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11709__A0 _11704_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12478_ _12472_/A _12478_/B vssd1 vssd1 vccd1 vccd1 _12479_/A sky130_fd_sc_hd__and2b_1
X_14217_ _13806_/X _14215_/B _14216_/Y _14000_/X vssd1 vssd1 vccd1 vccd1 _14217_/X
+ sky130_fd_sc_hd__o211a_1
X_17005_ _17062_/S vssd1 vssd1 vccd1 vccd1 _17014_/S sky130_fd_sc_hd__buf_2
X_11429_ _18300_/Q vssd1 vssd1 vccd1 vccd1 _12765_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15197_ _16699_/A vssd1 vssd1 vccd1 vccd1 _15197_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14148_ _12066_/Y _14070_/X _14147_/X _14099_/X vssd1 vssd1 vccd1 vccd1 _14148_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17047__S _17047_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11884__A _19667_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18956_ _19414_/CLK _18956_/D vssd1 vssd1 vccd1 vccd1 _18956_/Q sky130_fd_sc_hd__dfxtp_1
X_14079_ _14075_/B _14074_/B _14077_/X _14078_/Y vssd1 vssd1 vccd1 vccd1 _14079_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17907_ _17909_/A _17907_/B vssd1 vssd1 vccd1 vccd1 _17908_/A sky130_fd_sc_hd__and2_1
XFILLER_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12685__A1 _18622_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18887_ _19442_/CLK _18887_/D vssd1 vssd1 vccd1 vccd1 _18887_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11032__S1 _10739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12685__B2 _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17073__A0 _16755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17838_ _15216_/X _19720_/Q _17838_/S vssd1 vssd1 vccd1 vccd1 _17839_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12437__A1 _19689_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17769_ _19689_/Q _17708_/A _17767_/Y _17768_/X vssd1 vssd1 vccd1 vccd1 _19689_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_81_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09302__A1 _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13604__A _13604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19508_ _19636_/CLK _19508_/D vssd1 vssd1 vccd1 vccd1 _19508_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09302__B2 _13523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19439_ _19601_/CLK _19439_/D vssd1 vssd1 vccd1 vccd1 _19439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17510__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_9_0_clock_A clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09123_ _18557_/Q _14511_/A _11297_/B _11297_/C vssd1 vssd1 vccd1 vccd1 _11343_/C
+ sky130_fd_sc_hd__and4bb_2
XANTENNA__16126__S _16129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11497__C _18563_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17300__A1 _16715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15266__A _16430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ _09874_/S _09954_/Y _09955_/Y _09881_/A vssd1 vssd1 vccd1 vccd1 _09956_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__14665__A2 _12660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12676__A1 _18335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09887_ _18842_/Q _19396_/Q _19558_/Q _18810_/Q _09809_/X _09881_/X vssd1 vssd1 vccd1
+ vccd1 _09888_/B sky130_fd_sc_hd__mux4_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15205__S _15217_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10800_ _19505_/Q _19119_/Q _19569_/Q _18725_/Q _10631_/A _10772_/X vssd1 vssd1 vccd1
+ vccd1 _10801_/B sky130_fd_sc_hd__mux4_2
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _11779_/Y _18495_/Q _11840_/A vssd1 vssd1 vccd1 vccd1 _13630_/A sky130_fd_sc_hd__mux2_4
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10857__B _10857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10731_ _09926_/A _10705_/Y _10730_/X _09305_/A _18433_/Q vssd1 vssd1 vccd1 vccd1
+ _10732_/A sky130_fd_sc_hd__a32o_4
XFILLER_159_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17420__S _17424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13450_ _13450_/A vssd1 vssd1 vccd1 vccd1 _18385_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13928__A1 _11602_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10662_ _10959_/A vssd1 vssd1 vccd1 vccd1 _10663_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__13928__B2 _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12401_ _12401_/A vssd1 vssd1 vccd1 vccd1 _14308_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_166_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13381_ _19686_/Q _13251_/X _12743_/X _18410_/Q vssd1 vssd1 vccd1 vccd1 _13381_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10873__A _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ _10593_/A _10593_/B vssd1 vssd1 vccd1 vccd1 _10593_/X sky130_fd_sc_hd__or2_1
XFILLER_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15120_ _18640_/Q _15116_/X _15118_/X _10051_/A vssd1 vssd1 vccd1 vccd1 _18640_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12332_ _12371_/A _12290_/B _12313_/A _12331_/X vssd1 vssd1 vccd1 vccd1 _12333_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_154_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09439__A _09629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15051_ _18455_/Q _13411_/B _15051_/S vssd1 vssd1 vccd1 vccd1 _15051_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12263_ _13615_/A vssd1 vssd1 vccd1 vccd1 _14227_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_108_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14002_ _14019_/S _14001_/Y _13706_/A vssd1 vssd1 vccd1 vccd1 _14002_/X sky130_fd_sc_hd__a21o_1
XFILLER_135_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11214_ _11365_/B vssd1 vssd1 vccd1 vccd1 _11282_/A sky130_fd_sc_hd__clkbuf_2
X_12194_ _11980_/X _12190_/X _12192_/X _12193_/X vssd1 vssd1 vccd1 vccd1 _12194_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18810_ _19590_/CLK _18810_/D vssd1 vssd1 vccd1 vccd1 _18810_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput73 _12511_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[0] sky130_fd_sc_hd__buf_2
X_11145_ _11145_/A vssd1 vssd1 vccd1 vccd1 _11145_/Y sky130_fd_sc_hd__inv_2
X_19790_ _19790_/CLK _19790_/D vssd1 vssd1 vccd1 vccd1 _19790_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput84 _11624_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[1] sky130_fd_sc_hd__buf_2
XANTENNA__10812__S _11028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput95 _11667_/B vssd1 vssd1 vccd1 vccd1 io_dbus_addr[2] sky130_fd_sc_hd__buf_2
XANTENNA__13313__C1 _13282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18741_ _19716_/CLK _18741_/D vssd1 vssd1 vccd1 vccd1 _18741_/Q sky130_fd_sc_hd__dfxtp_1
X_15953_ _17892_/A vssd1 vssd1 vccd1 vccd1 _17779_/A sky130_fd_sc_hd__clkbuf_1
X_11076_ _10881_/X _11073_/X _11257_/B _11254_/C _11252_/A vssd1 vssd1 vccd1 vccd1
+ _11248_/B sky130_fd_sc_hd__a2111o_1
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10027_ _10007_/X _10020_/X _10022_/X _10026_/X _09249_/A vssd1 vssd1 vccd1 vccd1
+ _10027_/X sky130_fd_sc_hd__a311o_1
XANTENNA__15904__A _15950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_1_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14904_ _14925_/A vssd1 vssd1 vccd1 vccd1 _14904_/X sky130_fd_sc_hd__buf_2
XANTENNA__17391__A _17391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18672_ _19295_/CLK _18672_/D vssd1 vssd1 vccd1 vccd1 _18672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15884_ _15884_/A vssd1 vssd1 vccd1 vccd1 _18945_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11082__A_N _12478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10773__S0 _10719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17623_ _17632_/C _17623_/B vssd1 vssd1 vccd1 vccd1 _17623_/Y sky130_fd_sc_hd__nand2_2
XFILLER_91_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14835_ _14833_/X _18596_/Q _14880_/S vssd1 vssd1 vccd1 vccd1 _14836_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13616__A0 _14045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17554_ _17554_/A vssd1 vssd1 vccd1 vccd1 _19636_/D sky130_fd_sc_hd__clkbuf_1
X_11978_ _11978_/A _11978_/B vssd1 vssd1 vccd1 vccd1 _11978_/X sky130_fd_sc_hd__xor2_4
X_14766_ _14766_/A _14786_/C vssd1 vssd1 vccd1 vccd1 _14766_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10525__S0 _10387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16505_ _16573_/S vssd1 vssd1 vccd1 vccd1 _16514_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_60_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10929_ _10996_/A _10926_/X _10928_/X _10821_/X vssd1 vssd1 vccd1 vccd1 _10929_/X
+ sky130_fd_sc_hd__o211a_1
X_13717_ _13785_/A _13720_/B _13720_/A vssd1 vssd1 vccd1 vccd1 _13974_/A sky130_fd_sc_hd__and3b_1
X_14697_ _14589_/A _14648_/X _14649_/X input58/X vssd1 vssd1 vccd1 vccd1 _14698_/B
+ sky130_fd_sc_hd__a22o_1
X_17485_ _19606_/Q _16670_/X _17485_/S vssd1 vssd1 vccd1 vccd1 _17486_/A sky130_fd_sc_hd__mux2_1
X_19224_ _19640_/CLK _19224_/D vssd1 vssd1 vccd1 vccd1 _19224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16436_ _16039_/X _19180_/Q _16442_/S vssd1 vssd1 vccd1 vccd1 _16437_/A sky130_fd_sc_hd__mux2_1
X_13648_ _13646_/X _13647_/X _13741_/S vssd1 vssd1 vccd1 vccd1 _13648_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ _19704_/CLK _19155_/D vssd1 vssd1 vccd1 vccd1 _19155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16367_ _19150_/Q _15500_/X _16369_/S vssd1 vssd1 vccd1 vccd1 _16368_/A sky130_fd_sc_hd__mux2_1
X_13579_ _13579_/A _13579_/B _13579_/C _13579_/D vssd1 vssd1 vccd1 vccd1 _13580_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18106_ _19822_/Q _18104_/B _18105_/Y vssd1 vssd1 vccd1 vccd1 _19822_/D sky130_fd_sc_hd__o21a_1
XFILLER_173_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15318_ _18711_/Q _15210_/X _15322_/S vssd1 vssd1 vccd1 vccd1 _15319_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19086_ _19568_/CLK _19086_/D vssd1 vssd1 vccd1 vccd1 _19086_/Q sky130_fd_sc_hd__dfxtp_1
X_16298_ _16355_/S vssd1 vssd1 vccd1 vccd1 _16307_/S sky130_fd_sc_hd__buf_2
XANTENNA__13147__A2 _13123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15785__S _15791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18037_ _18071_/A _18043_/C vssd1 vssd1 vccd1 vccd1 _18037_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_79_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15249_ _18684_/Q _15248_/X _15260_/S vssd1 vssd1 vccd1 vccd1 _15250_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11158__A1 _09172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09810_ _09810_/A vssd1 vssd1 vccd1 vccd1 _09810_/X sky130_fd_sc_hd__buf_2
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12503__A _12503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09741_ _09318_/A _09725_/Y _09731_/X _09740_/Y _09395_/A vssd1 vssd1 vccd1 vccd1
+ _09741_/X sky130_fd_sc_hd__o311a_2
X_18939_ _19722_/CLK _18939_/D vssd1 vssd1 vccd1 vccd1 _18939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11119__A _11119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17505__S _17507_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ _10401_/A vssd1 vssd1 vccd1 vccd1 _09673_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_67_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11553__S _14032_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10436__A3 _10435_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14032__A0 _18434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14583__A1 _11517_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10819__S1 _10739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09106_ _09119_/A vssd1 vssd1 vccd1 vccd1 _09106_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_109_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17476__A _17533_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09939_ _09879_/A _09934_/X _09938_/X _09320_/A vssd1 vssd1 vccd1 vccd1 _09940_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13228__B _13228_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12950_ _18293_/Q _12952_/C _12949_/Y vssd1 vssd1 vccd1 vccd1 _18293_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__13310__A2 _13307_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17588__A1 _16819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ _11901_/A _19737_/Q _11901_/C vssd1 vssd1 vccd1 vccd1 _11984_/D sky130_fd_sc_hd__and3_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09722__A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12881_ _12883_/B _12883_/C _12880_/Y vssd1 vssd1 vccd1 vccd1 _18273_/D sky130_fd_sc_hd__o21a_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13244__A _18628_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _14624_/A _14620_/B vssd1 vssd1 vccd1 vccd1 _14621_/A sky130_fd_sc_hd__and2_1
X_11832_ _11911_/C vssd1 vssd1 vccd1 vccd1 _12023_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14551_/A _14551_/B vssd1 vssd1 vccd1 vccd1 _14551_/Y sky130_fd_sc_hd__nand2_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _18349_/Q _18382_/Q _11720_/B _11762_/X vssd1 vssd1 vccd1 vccd1 _11764_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14774__S _14822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _18409_/Q _13376_/X _13508_/S vssd1 vssd1 vccd1 vccd1 _13503_/A sky130_fd_sc_hd__mux2_1
X_10714_ _10788_/S _10666_/Y _10711_/Y _10713_/X vssd1 vssd1 vccd1 vccd1 _10714_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10832__B1 _10821_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ _17270_/A vssd1 vssd1 vccd1 vccd1 _19510_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _14482_/A vssd1 vssd1 vccd1 vccd1 _18511_/D sky130_fd_sc_hd__clkbuf_1
X_11694_ _12463_/A _11693_/X _11835_/S vssd1 vssd1 vccd1 vccd1 _13653_/A sky130_fd_sc_hd__mux2_4
XANTENNA__17760__A1 _19687_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13433_ _18266_/Q _12582_/X _12584_/X _19855_/Q _13432_/X vssd1 vssd1 vccd1 vccd1
+ _13433_/X sky130_fd_sc_hd__a221o_1
X_16221_ _16221_/A vssd1 vssd1 vccd1 vccd1 _19085_/D sky130_fd_sc_hd__clkbuf_1
X_10645_ _10764_/A _10645_/B vssd1 vssd1 vccd1 vccd1 _10645_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16152_ _16209_/S vssd1 vssd1 vccd1 vccd1 _16161_/S sky130_fd_sc_hd__buf_2
X_13364_ _12577_/X _13355_/Y _13363_/X _12596_/X _18644_/Q vssd1 vssd1 vccd1 vccd1
+ _13364_/X sky130_fd_sc_hd__a32o_4
XANTENNA__09169__A _09169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10576_ _10475_/A _10575_/X _09459_/A vssd1 vssd1 vccd1 vccd1 _10576_/X sky130_fd_sc_hd__o21a_1
XFILLER_155_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12315_ _12315_/A _12335_/C vssd1 vssd1 vccd1 vccd1 _12315_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_80_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15103_ _18628_/Q _15102_/X _15097_/X _10601_/B vssd1 vssd1 vccd1 vccd1 _18628_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16083_ _16793_/A vssd1 vssd1 vccd1 vccd1 _16083_/X sky130_fd_sc_hd__clkbuf_1
X_13295_ _13295_/A _13295_/B vssd1 vssd1 vccd1 vccd1 _13295_/X sky130_fd_sc_hd__or2_1
XANTENNA__12337__A0 _12333_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14803__A _14842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15034_ _15033_/X _18613_/Q _15056_/S vssd1 vssd1 vccd1 vccd1 _15035_/A sky130_fd_sc_hd__mux2_1
X_12246_ _12246_/A _12267_/C vssd1 vssd1 vccd1 vccd1 _12246_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19842_ _19851_/CLK _19842_/D vssd1 vssd1 vccd1 vccd1 _19842_/Q sky130_fd_sc_hd__dfxtp_1
X_12177_ _12177_/A vssd1 vssd1 vccd1 vccd1 _12444_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_111_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ _09428_/A _11117_/X _11126_/X _09625_/A _11127_/Y vssd1 vssd1 vccd1 vccd1
+ _12481_/A sky130_fd_sc_hd__o32a_4
X_19773_ _19779_/CLK _19773_/D vssd1 vssd1 vccd1 vccd1 _19773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16985_ _16985_/A vssd1 vssd1 vccd1 vccd1 _19399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18724_ _19632_/CLK _18724_/D vssd1 vssd1 vccd1 vccd1 _18724_/Q sky130_fd_sc_hd__dfxtp_1
X_15936_ _15936_/A vssd1 vssd1 vccd1 vccd1 _18969_/D sky130_fd_sc_hd__clkbuf_1
X_11059_ _19501_/Q _19115_/Q _19565_/Q _18721_/Q _10710_/A _09480_/A vssd1 vssd1 vccd1
+ vccd1 _11060_/B sky130_fd_sc_hd__mux4_2
XFILLER_77_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09632__A _09632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18655_ _19700_/CLK _18655_/D vssd1 vssd1 vccd1 vccd1 _18655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15867_ _15867_/A vssd1 vssd1 vccd1 vccd1 _18938_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10778__A _10807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17606_ _17606_/A vssd1 vssd1 vccd1 vccd1 _19660_/D sky130_fd_sc_hd__clkbuf_1
X_14818_ input32/X _14801_/X _14804_/X vssd1 vssd1 vccd1 vccd1 _14818_/X sky130_fd_sc_hd__a21o_1
X_18586_ _19696_/CLK _18586_/D vssd1 vssd1 vccd1 vccd1 _18586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15798_ _15033_/X _18908_/Q _15802_/S vssd1 vssd1 vccd1 vccd1 _15799_/A sky130_fd_sc_hd__mux2_1
X_17537_ _17605_/S vssd1 vssd1 vccd1 vccd1 _17546_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_33_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14749_ _14981_/S _12683_/B _14747_/Y _14945_/B vssd1 vssd1 vccd1 vccd1 _14749_/X
+ sky130_fd_sc_hd__a211o_2
XANTENNA__17060__S _17062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17468_ _19598_/Q _16645_/X _17474_/S vssd1 vssd1 vccd1 vccd1 _17469_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19207_ _19271_/CLK _19207_/D vssd1 vssd1 vccd1 vccd1 _19207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16419_ _16419_/A vssd1 vssd1 vccd1 vccd1 _19173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_182_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19541_/CLK sky130_fd_sc_hd__clkbuf_16
X_17399_ _17399_/A vssd1 vssd1 vccd1 vccd1 _19567_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09667__S1 _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19138_ _19427_/CLK _19138_/D vssd1 vssd1 vccd1 vccd1 _19138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14317__A1 _12408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19069_ _19718_/CLK _19069_/D vssd1 vssd1 vccd1 vccd1 _19069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_120_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _18548_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09724_ _19269_/Q _19040_/Q _18971_/Q _19365_/Q _09721_/X _09723_/X vssd1 vssd1 vccd1
+ vccd1 _09725_/B sky130_fd_sc_hd__mux4_1
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09542__A _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ _09649_/A _09652_/X _09654_/X _09708_/A vssd1 vssd1 vccd1 vccd1 _09655_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_135_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19693_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09586_ _10331_/A _09585_/X vssd1 vssd1 vccd1 vccd1 _09586_/X sky130_fd_sc_hd__or2b_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10290__A1 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_102_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10430_ _10432_/A _10429_/X _09212_/A vssd1 vssd1 vccd1 vccd1 _10430_/X sky130_fd_sc_hd__o21a_1
XFILLER_164_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10361_ _10477_/A vssd1 vssd1 vccd1 vccd1 _10428_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16314__S _16318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12319__B1 _18375_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12100_ _13312_/A _12123_/C _17241_/S vssd1 vssd1 vccd1 vccd1 _12100_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13080_ _18341_/Q _12564_/A _12585_/A _18274_/Q _12640_/A vssd1 vssd1 vccd1 vccd1
+ _13080_/X sky130_fd_sc_hd__a221o_1
XANTENNA__09717__A _10262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10292_ _11123_/A _10292_/B vssd1 vssd1 vccd1 vccd1 _10292_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12031_ _12057_/A _12131_/B vssd1 vssd1 vccd1 vccd1 _12032_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13531__A2 _12692_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_1_1_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14769__S _14923_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16770_ _16770_/A vssd1 vssd1 vccd1 vccd1 _19314_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14492__A0 _18516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13982_ _14003_/A vssd1 vssd1 vccd1 vccd1 _13982_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15721_ _15721_/A vssd1 vssd1 vccd1 vccd1 _15730_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12933_ _18288_/Q _18287_/Q _12933_/C _12933_/D vssd1 vssd1 vccd1 vccd1 _12934_/A
+ sky130_fd_sc_hd__and4_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_27_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16984__S _16986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _19695_/CLK _18440_/D vssd1 vssd1 vccd1 vccd1 _18440_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _18843_/Q _15574_/X _15658_/S vssd1 vssd1 vccd1 vccd1 _15653_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12864_ _12904_/A _12864_/B _12864_/C vssd1 vssd1 vccd1 vccd1 _18268_/D sky130_fd_sc_hd__nor3_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14603_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18371_ _19082_/CLK _18371_/D vssd1 vssd1 vccd1 vccd1 _18371_/Q sky130_fd_sc_hd__dfxtp_2
X_11815_ _11849_/A _12095_/B vssd1 vssd1 vccd1 vccd1 _11815_/X sky130_fd_sc_hd__xor2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12795_ _19860_/Q _19859_/Q _18214_/B _18214_/C vssd1 vssd1 vccd1 vccd1 _18222_/C
+ sky130_fd_sc_hd__and4_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output101_A _11813_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _16838_/A vssd1 vssd1 vccd1 vccd1 _15583_/X sky130_fd_sc_hd__buf_2
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16285__A _17391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13702__A _13702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17322_ _16743_/X _19533_/Q _17330_/S vssd1 vssd1 vccd1 vccd1 _17323_/A sky130_fd_sc_hd__mux2_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14534_ _17892_/A vssd1 vssd1 vccd1 vccd1 _14585_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11746_ _11746_/A _11746_/B vssd1 vssd1 vccd1 vccd1 _11747_/B sky130_fd_sc_hd__nor2_2
XFILLER_30_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10900__S0 _10724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10281__A1 _09735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17253_ _17253_/A vssd1 vssd1 vccd1 vccd1 _19502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11677_ _18350_/Q _15263_/A vssd1 vssd1 vccd1 vccd1 _11827_/B sky130_fd_sc_hd__nand2_2
X_14465_ _18504_/Q _12067_/B _14465_/S vssd1 vssd1 vccd1 vccd1 _14466_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16204_ _16204_/A vssd1 vssd1 vccd1 vccd1 _19074_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11222__A _11222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13416_ _18297_/Q _12606_/A _12546_/A _18380_/Q _12641_/A vssd1 vssd1 vccd1 vccd1
+ _13416_/X sky130_fd_sc_hd__a221o_1
X_10628_ _09451_/A _10625_/X _10627_/X _09225_/A vssd1 vssd1 vccd1 vccd1 _10628_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09423__B1 _09415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17184_ _18439_/Q _13279_/X _17184_/S vssd1 vssd1 vccd1 vccd1 _17184_/X sky130_fd_sc_hd__mux2_1
X_14396_ _14396_/A vssd1 vssd1 vccd1 vccd1 _18477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13347_ _18372_/Q _13352_/B vssd1 vssd1 vccd1 vccd1 _13347_/X sky130_fd_sc_hd__or2_1
X_16135_ _16134_/X _19045_/Q _16135_/S vssd1 vssd1 vccd1 vccd1 _16136_/A sky130_fd_sc_hd__mux2_1
X_10559_ _10559_/A _10559_/B vssd1 vssd1 vccd1 vccd1 _10559_/X sky130_fd_sc_hd__and2_1
XFILLER_143_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14533__A _18563_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16224__S _16224_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13278_ _18632_/Q _14859_/B _14859_/C _14859_/D vssd1 vssd1 vccd1 vccd1 _13278_/X
+ sky130_fd_sc_hd__or4_1
X_16066_ _16066_/A vssd1 vssd1 vccd1 vccd1 _19023_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12229_ _12106_/A _14216_/A _12205_/B vssd1 vssd1 vccd1 vccd1 _12230_/B sky130_fd_sc_hd__o21a_1
X_15017_ _18452_/Q _14958_/A _14829_/B vssd1 vssd1 vccd1 vccd1 _15017_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_111_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19825_ _19866_/CLK _19825_/D vssd1 vssd1 vccd1 vccd1 _19825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15364__A _15410_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19756_ _19759_/CLK _19756_/D vssd1 vssd1 vccd1 vccd1 _19756_/Q sky130_fd_sc_hd__dfxtp_4
X_16968_ _16968_/A vssd1 vssd1 vccd1 vccd1 _19391_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_52_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19427_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13286__B2 _13295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__A _09810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18707_ _19645_/CLK _18707_/D vssd1 vssd1 vccd1 vccd1 _18707_/Q sky130_fd_sc_hd__dfxtp_1
X_15919_ _15919_/A vssd1 vssd1 vccd1 vccd1 _18961_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16894__S _16902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19687_ _19687_/CLK _19687_/D vssd1 vssd1 vccd1 vccd1 _19687_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16899_ _16899_/A vssd1 vssd1 vccd1 vccd1 _19361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09440_ _10540_/S vssd1 vssd1 vccd1 vccd1 _10350_/S sky130_fd_sc_hd__buf_4
XFILLER_80_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14235__A0 _18448_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18638_ _19081_/CLK _18638_/D vssd1 vssd1 vccd1 vccd1 _18638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09371_ _09370_/A _09368_/Y _09370_/Y _09421_/A vssd1 vssd1 vccd1 vccd1 _09371_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18569_ _18578_/CLK _18569_/D vssd1 vssd1 vccd1 vccd1 _18569_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_67_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _18330_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15303__S _15311_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11772__B2 _11788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09537__A _10262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17660__A0 _19669_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13277__A1 _19837_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09272__A _10857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09707_ _10262_/A _09707_/B vssd1 vssd1 vccd1 vccd1 _09707_/X sky130_fd_sc_hd__or2_1
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11288__B1 _11278_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09638_ _10309_/A _09638_/B vssd1 vssd1 vccd1 vccd1 _09638_/X sky130_fd_sc_hd__or2_1
XFILLER_71_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14777__A1 _13211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09569_ _18846_/Q _19400_/Q _19562_/Q _18814_/Q _09553_/X _09555_/X vssd1 vssd1 vccd1
+ vccd1 _09569_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14618__A _14638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11600_ _11534_/A _13526_/C _11565_/C _11287_/X vssd1 vssd1 vccd1 vccd1 _13572_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12580_ _18252_/Q vssd1 vssd1 vccd1 vccd1 _12808_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17715__A1 _19678_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10263__A1 _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11531_ _11531_/A _11640_/A _11640_/B vssd1 vssd1 vccd1 vccd1 _11531_/X sky130_fd_sc_hd__or3_1
XFILLER_157_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14250_ _14250_/A _14253_/A vssd1 vssd1 vccd1 vccd1 _14250_/Y sky130_fd_sc_hd__nor2_1
X_11462_ _11462_/A _13532_/A vssd1 vssd1 vccd1 vccd1 _12658_/A sky130_fd_sc_hd__or2_4
XFILLER_165_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13201_ _13185_/X _13197_/X _13200_/X _13167_/X vssd1 vssd1 vccd1 vccd1 _18355_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_137_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09956__A1 _09874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10413_ _10413_/A _10413_/B vssd1 vssd1 vccd1 vccd1 _10414_/A sky130_fd_sc_hd__or2_1
XFILLER_125_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14181_ _14178_/B _14176_/B _13721_/X _14179_/X _14180_/X vssd1 vssd1 vccd1 vccd1
+ _14182_/B sky130_fd_sc_hd__o221a_1
XFILLER_165_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11393_ _18549_/Q _18548_/Q _18547_/Q _18546_/Q vssd1 vssd1 vccd1 vccd1 _11412_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_165_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13132_ _18303_/Q _13130_/X _12665_/A _19792_/Q _13131_/X vssd1 vssd1 vccd1 vccd1
+ _13132_/X sky130_fd_sc_hd__a221o_1
XFILLER_48_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input62_A io_ibus_inst[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09447__A _09447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ _10337_/Y _10339_/Y _10341_/Y _10343_/Y _09403_/A vssd1 vssd1 vccd1 vccd1
+ _10344_/X sky130_fd_sc_hd__o221a_2
XFILLER_140_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11188__S _11188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15883__S _15891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17940_ _17944_/B _17944_/C _13063_/X vssd1 vssd1 vccd1 vccd1 _17940_/Y sky130_fd_sc_hd__a21oi_1
X_13063_ _17993_/A vssd1 vssd1 vccd1 vccd1 _13063_/X sky130_fd_sc_hd__clkbuf_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10275_ _19259_/Q _19030_/Q _18961_/Q _19355_/Q _09675_/S _10239_/X vssd1 vssd1 vccd1
+ vccd1 _10276_/B sky130_fd_sc_hd__mux4_1
XFILLER_140_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10949__S0 _10719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ _19741_/Q vssd1 vssd1 vccd1 vccd1 _12043_/A sky130_fd_sc_hd__buf_4
XFILLER_105_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17871_ _17871_/A vssd1 vssd1 vccd1 vccd1 _19736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19610_ _19610_/CLK _19610_/D vssd1 vssd1 vccd1 vccd1 _19610_/Q sky130_fd_sc_hd__dfxtp_1
X_16822_ _16822_/A vssd1 vssd1 vccd1 vccd1 _16822_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15184__A _16686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14465__A0 _18504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09182__A _11099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09567__S0 _09553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19541_ _19541_/CLK _19541_/D vssd1 vssd1 vccd1 vccd1 _19541_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11279__B1 _11278_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16753_ _16752_/X _19309_/Q _16759_/S vssd1 vssd1 vccd1 vccd1 _16754_/A sky130_fd_sc_hd__mux2_1
X_13965_ _13839_/X _13964_/Y _13965_/S vssd1 vssd1 vccd1 vccd1 _13965_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17603__S _17605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15704_ _18866_/Q _15545_/X _15708_/S vssd1 vssd1 vccd1 vccd1 _15705_/A sky130_fd_sc_hd__mux2_1
X_12916_ _12925_/C _12919_/C _12915_/Y vssd1 vssd1 vccd1 vccd1 _18283_/D sky130_fd_sc_hd__o21a_1
X_19472_ _19472_/CLK _19472_/D vssd1 vssd1 vccd1 vccd1 _19472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16684_ _19288_/Q _16683_/X _16687_/S vssd1 vssd1 vccd1 vccd1 _16685_/A sky130_fd_sc_hd__mux2_1
X_13896_ _14182_/A vssd1 vssd1 vccd1 vccd1 _14130_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10510__A_N _10384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18423_ _19468_/CLK _18423_/D vssd1 vssd1 vccd1 vccd1 _18423_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__14768__A1 _13196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15635_ _15635_/A vssd1 vssd1 vccd1 vccd1 _18835_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _12850_/B _12850_/C _12817_/X vssd1 vssd1 vccd1 vccd1 _12847_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _18386_/CLK _18354_/D vssd1 vssd1 vccd1 vccd1 _18354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15566_ _15566_/A vssd1 vssd1 vccd1 vccd1 _18808_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _18643_/Q _12778_/B vssd1 vssd1 vccd1 vccd1 _12778_/X sky130_fd_sc_hd__or2_1
XFILLER_30_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17305_ _19526_/Q _16721_/X _17313_/S vssd1 vssd1 vccd1 vccd1 _17306_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14517_ _17862_/A _14517_/B vssd1 vssd1 vccd1 vccd1 _14518_/A sky130_fd_sc_hd__or2_1
XFILLER_30_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18285_ _19759_/CLK _18285_/D vssd1 vssd1 vccd1 vccd1 _18285_/Q sky130_fd_sc_hd__dfxtp_1
X_11729_ _11729_/A vssd1 vssd1 vccd1 vccd1 _11801_/A sky130_fd_sc_hd__clkbuf_2
X_15497_ _16752_/A vssd1 vssd1 vccd1 vccd1 _15497_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17236_ _19497_/Q _17235_/X _17239_/S vssd1 vssd1 vccd1 vccd1 _17237_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14448_ _18496_/Q _11849_/A _14454_/S vssd1 vssd1 vccd1 vccd1 _14449_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17167_ _18434_/Q _13230_/X _17167_/S vssd1 vssd1 vccd1 vccd1 _17167_/X sky130_fd_sc_hd__mux2_1
X_14379_ _14379_/A vssd1 vssd1 vccd1 vccd1 _18471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12951__B1 _18294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16118_ _16118_/A vssd1 vssd1 vccd1 vccd1 _19039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09357__A _11113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17098_ _17098_/A vssd1 vssd1 vccd1 vccd1 _19449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16889__S _16891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16049_ _16048_/X _19018_/Q _16049_/S vssd1 vssd1 vccd1 vccd1 _16050_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10714__C1 _10713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15248__A2 _13136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17642__A0 _13088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19808_ _19810_/CLK _19808_/D vssd1 vssd1 vccd1 vccd1 _19808_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13607__A _13607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13259__B2 _18629_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10190__B1 _09317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19739_ _19753_/CLK _19739_/D vssd1 vssd1 vccd1 vccd1 _19739_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__10168__S1 _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11127__A _18439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09423_ _09814_/A _09422_/X _09415_/X vssd1 vssd1 vccd1 vccd1 _09423_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_92_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14759__A1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14759__B2 _14732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16129__S _16129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09354_ _10651_/A vssd1 vssd1 vccd1 vccd1 _10384_/A sky130_fd_sc_hd__buf_2
XFILLER_12_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13431__B2 _19690_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15968__S _15972_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09285_ _09285_/A vssd1 vssd1 vccd1 vccd1 _09285_/X sky130_fd_sc_hd__buf_2
XFILLER_139_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15269__A _15337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10905__S _10905_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10953__C1 _09391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10206__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09797__S0 _09976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10060_ _19423_/Q _19199_/Q _19716_/Q _19167_/Q _09808_/A _09936_/A vssd1 vssd1 vccd1
+ vccd1 _10060_/X sky130_fd_sc_hd__mux4_1
XFILLER_134_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15208__S _15217_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13517__A _13563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18189__A1 _19850_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13750_ _13969_/S vssd1 vssd1 vccd1 vccd1 _13750_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10962_ _10992_/A _10962_/B vssd1 vssd1 vccd1 vccd1 _10962_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13670__A1 _12510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12701_ _13426_/A _18630_/Q vssd1 vssd1 vccd1 vccd1 _12701_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09730__A _09867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13681_ _12262_/B _14026_/B _13681_/S vssd1 vssd1 vccd1 vccd1 _13681_/X sky130_fd_sc_hd__mux2_1
X_10893_ _10793_/X _10883_/Y _10888_/X _10892_/Y _09391_/A vssd1 vssd1 vccd1 vccd1
+ _10893_/X sky130_fd_sc_hd__o311a_1
XANTENNA__11108__S0 _10279_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15420_ _18754_/Q _15143_/X _15426_/S vssd1 vssd1 vccd1 vccd1 _15421_/A sky130_fd_sc_hd__mux2_1
X_12632_ _18638_/Q _12632_/B vssd1 vssd1 vccd1 vccd1 _12632_/X sky130_fd_sc_hd__or2_1
XFILLER_169_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15878__S _15878_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12563_ _12563_/A vssd1 vssd1 vccd1 vccd1 _12564_/A sky130_fd_sc_hd__clkbuf_2
X_15351_ _18725_/Q _15152_/X _15351_/S vssd1 vssd1 vccd1 vccd1 _15352_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14302_ _13788_/A _14299_/X _14301_/Y _13894_/A vssd1 vssd1 vccd1 vccd1 _14302_/X
+ sky130_fd_sc_hd__a31o_1
X_11514_ _11514_/A vssd1 vssd1 vccd1 vccd1 _11517_/B sky130_fd_sc_hd__clkbuf_4
X_18070_ _18070_/A vssd1 vssd1 vccd1 vccd1 _18075_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15282_ _15282_/A vssd1 vssd1 vccd1 vccd1 _18694_/D sky130_fd_sc_hd__clkbuf_1
X_12494_ _12494_/A vssd1 vssd1 vccd1 vccd1 _12494_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09929__A1 _09928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17021_ _19415_/Q _16680_/X _17025_/S vssd1 vssd1 vccd1 vccd1 _17022_/A sky130_fd_sc_hd__mux2_1
X_11445_ _18346_/Q _18339_/Q _18340_/Q _18347_/Q vssd1 vssd1 vccd1 vccd1 _11721_/A
+ sky130_fd_sc_hd__a22o_1
X_14233_ _14426_/A vssd1 vssd1 vccd1 vccd1 _14384_/A sky130_fd_sc_hd__buf_2
XANTENNA__14922__A1 _12615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14164_ _14168_/A _14168_/B vssd1 vssd1 vccd1 vccd1 _14164_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09177__A _09177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11376_ _11376_/A _11534_/B _11376_/C _11322_/D vssd1 vssd1 vccd1 vccd1 _11531_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13115_ _13115_/A vssd1 vssd1 vccd1 vccd1 _13119_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10327_ _10327_/A _10327_/B vssd1 vssd1 vccd1 vccd1 _10327_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14095_ _13862_/A _14090_/X _14092_/Y _14094_/X vssd1 vssd1 vccd1 vccd1 _14095_/X
+ sky130_fd_sc_hd__o31a_1
X_18972_ _19723_/CLK _18972_/D vssd1 vssd1 vccd1 vccd1 _18972_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13489__A1 _12656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17923_ _17927_/D vssd1 vssd1 vccd1 vccd1 _18105_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13046_ _17935_/A _13046_/B _13046_/C vssd1 vssd1 vccd1 vccd1 _18326_/D sky130_fd_sc_hd__nor3_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10258_ _09173_/A _10257_/X _09772_/A vssd1 vssd1 vccd1 vccd1 _10258_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17624__A0 _13182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09624__B _09624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17854_ _17854_/A vssd1 vssd1 vccd1 vccd1 _19727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10189_ _19421_/Q _19197_/Q _19714_/Q _19165_/Q _10129_/S _09723_/A vssd1 vssd1 vccd1
+ vccd1 _10189_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16805_ _16805_/A vssd1 vssd1 vccd1 vccd1 _19325_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14646__A1_N input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14989__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17785_ _17853_/S vssd1 vssd1 vccd1 vccd1 _17794_/S sky130_fd_sc_hd__clkbuf_4
X_14997_ _14996_/X _18610_/Q _14997_/S vssd1 vssd1 vccd1 vccd1 _14998_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19524_ _19718_/CLK _19524_/D vssd1 vssd1 vccd1 vccd1 _19524_/Q sky130_fd_sc_hd__dfxtp_1
X_16736_ _16736_/A vssd1 vssd1 vccd1 vccd1 _19304_/D sky130_fd_sc_hd__clkbuf_1
X_13948_ _13970_/S _13947_/X _13899_/X vssd1 vssd1 vccd1 vccd1 _13949_/B sky130_fd_sc_hd__o21ai_2
XFILLER_34_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09640__A _09640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19455_ _19716_/CLK _19455_/D vssd1 vssd1 vccd1 vccd1 _19455_/Q sky130_fd_sc_hd__dfxtp_1
X_16667_ _16667_/A vssd1 vssd1 vccd1 vccd1 _16667_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13879_ _13754_/X _13758_/X _13879_/S vssd1 vssd1 vccd1 vccd1 _13879_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18406_ _19788_/CLK _18406_/D vssd1 vssd1 vccd1 vccd1 _18406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15618_ _15618_/A vssd1 vssd1 vccd1 vccd1 _18827_/D sky130_fd_sc_hd__clkbuf_1
X_19386_ _19549_/CLK _19386_/D vssd1 vssd1 vccd1 vccd1 _19386_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09617__B1 _09616_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16598_ _16598_/A vssd1 vssd1 vccd1 vccd1 _19254_/D sky130_fd_sc_hd__clkbuf_1
X_18337_ _18401_/CLK _18337_/D vssd1 vssd1 vccd1 vccd1 _18337_/Q sky130_fd_sc_hd__dfxtp_1
X_15549_ _18803_/Q _15548_/X _15552_/S vssd1 vssd1 vccd1 vccd1 _15550_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15166__A1 _15165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18268_ _19472_/CLK _18268_/D vssd1 vssd1 vccd1 vccd1 _18268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17219_ _19492_/Q _17218_/X _17223_/S vssd1 vssd1 vccd1 vccd1 _17220_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_149_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18199_ _18199_/A vssd1 vssd1 vccd1 vccd1 _18223_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16920__B _16920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09972_ _09965_/X _09967_/X _09969_/X _09971_/X _09395_/X vssd1 vssd1 vccd1 vccd1
+ _09972_/X sky130_fd_sc_hd__a221o_2
XFILLER_131_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17615__A0 _19661_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09534__B _12504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14429__A0 _18489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09550__A _10475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14168__A _14168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09406_ _10774_/A vssd1 vssd1 vccd1 vccd1 _09407_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10218__B2 _18443_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09337_ _10706_/S vssd1 vssd1 vccd1 vccd1 _10836_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_138_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13800__A _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15157__A1 _15155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ _18573_/Q _18533_/Q vssd1 vssd1 vccd1 vccd1 _09268_/Y sky130_fd_sc_hd__xnor2_1
X_09199_ _09640_/A vssd1 vssd1 vccd1 vccd1 _11171_/A sky130_fd_sc_hd__buf_2
XFILLER_135_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12915__B1 _12869_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11230_ _11230_/A _11234_/A _11230_/C vssd1 vssd1 vccd1 vccd1 _11233_/A sky130_fd_sc_hd__and3_1
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ _18781_/Q _19010_/Q _18941_/Q _19239_/Q _09692_/A _10306_/A vssd1 vssd1 vccd1
+ vccd1 _11162_/B sky130_fd_sc_hd__mux4_1
XFILLER_106_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17418__S _17424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14631__A _14654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10112_ _10007_/X _10105_/X _10107_/X _10111_/X _09249_/A vssd1 vssd1 vccd1 vccd1
+ _10112_/X sky130_fd_sc_hd__a311o_1
XANTENNA__09725__A _10177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11092_ _18766_/Q _18995_/Q _18926_/Q _19224_/Q _09449_/A _09538_/A vssd1 vssd1 vccd1
+ vccd1 _11093_/B sky130_fd_sc_hd__mux4_1
XFILLER_121_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12143__A1 _19745_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13340__B1 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17942__A _18085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ _19650_/Q _19067_/Q _19104_/Q _18710_/Q _09952_/S _10029_/X vssd1 vssd1 vccd1
+ vccd1 _10044_/B sky130_fd_sc_hd__mux4_1
XFILLER_1_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14920_ _14920_/A vssd1 vssd1 vccd1 vccd1 _18603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input25_A io_dbus_rdata[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14851_ _14861_/A _14861_/C vssd1 vssd1 vccd1 vccd1 _14851_/X sky130_fd_sc_hd__xor2_1
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15093__A0 _18623_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13802_ _14040_/A vssd1 vssd1 vccd1 vccd1 _14088_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17570_ _17592_/A vssd1 vssd1 vccd1 vccd1 _17579_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_29_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14782_ _16765_/A vssd1 vssd1 vccd1 vccd1 _14782_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11994_ _11994_/A vssd1 vssd1 vccd1 vccd1 _12091_/A sky130_fd_sc_hd__clkbuf_2
X_16521_ _19218_/Q _15513_/X _16525_/S vssd1 vssd1 vccd1 vccd1 _16522_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10457__A1 _09681_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13733_ _13870_/A vssd1 vssd1 vccd1 vccd1 _13933_/A sky130_fd_sc_hd__clkbuf_2
X_10945_ _19504_/Q _19118_/Q _19568_/Q _18724_/Q _10706_/S _09481_/A vssd1 vssd1 vccd1
+ vccd1 _10946_/B sky130_fd_sc_hd__mux4_2
XFILLER_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19240_ _19725_/CLK _19240_/D vssd1 vssd1 vccd1 vccd1 _19240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16452_ _16452_/A vssd1 vssd1 vccd1 vccd1 _19187_/D sky130_fd_sc_hd__clkbuf_1
X_13664_ _13833_/B _13663_/X _13743_/S vssd1 vssd1 vccd1 vccd1 _13664_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10876_ _19634_/Q _19051_/Q _19088_/Q _18694_/Q _10614_/X _10616_/X vssd1 vssd1 vccd1
+ vccd1 _10876_/X sky130_fd_sc_hd__mux4_2
X_15403_ _15403_/A vssd1 vssd1 vccd1 vccd1 _18748_/D sky130_fd_sc_hd__clkbuf_1
X_19171_ _19557_/CLK _19171_/D vssd1 vssd1 vccd1 vccd1 _19171_/Q sky130_fd_sc_hd__dfxtp_1
X_12615_ _18637_/Q _12615_/B vssd1 vssd1 vccd1 vccd1 _12615_/X sky130_fd_sc_hd__or2_1
XFILLER_169_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16383_ _19157_/Q _15522_/X _16391_/S vssd1 vssd1 vccd1 vccd1 _16384_/A sky130_fd_sc_hd__mux2_1
X_13595_ _13595_/A vssd1 vssd1 vccd1 vccd1 _14111_/A sky130_fd_sc_hd__buf_2
XFILLER_129_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10304__S1 _09555_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18122_ _19828_/Q _19827_/Q _19826_/Q _18122_/D vssd1 vssd1 vccd1 vccd1 _18133_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_61_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15334_ _15334_/A vssd1 vssd1 vccd1 vccd1 _18718_/D sky130_fd_sc_hd__clkbuf_1
X_12546_ _12546_/A vssd1 vssd1 vccd1 vccd1 _12642_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18053_ _18077_/A _18053_/B _18053_/C vssd1 vssd1 vccd1 vccd1 _19803_/D sky130_fd_sc_hd__nor3_1
XANTENNA_clkbuf_leaf_150_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15265_ _15265_/A vssd1 vssd1 vccd1 vccd1 _18688_/D sky130_fd_sc_hd__clkbuf_1
X_12477_ _12477_/A vssd1 vssd1 vccd1 vccd1 _12477_/X sky130_fd_sc_hd__clkbuf_1
X_17004_ _17004_/A vssd1 vssd1 vccd1 vccd1 _19407_/D sky130_fd_sc_hd__clkbuf_1
X_14216_ _14216_/A _14216_/B vssd1 vssd1 vccd1 vccd1 _14216_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_output93_A _12385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11428_ _18551_/Q vssd1 vssd1 vccd1 vccd1 _11428_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15196_ _15196_/A vssd1 vssd1 vccd1 vccd1 _18668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14147_ _14054_/X _14137_/Y _14146_/X _14097_/X vssd1 vssd1 vccd1 vccd1 _14147_/X
+ sky130_fd_sc_hd__o211a_1
X_11359_ _11355_/Y _11343_/X _11356_/Y _11357_/Y _11584_/A vssd1 vssd1 vccd1 vccd1
+ _11587_/B sky130_fd_sc_hd__a32o_1
XFILLER_141_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14541__A _16430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09635__A _09635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18955_ _19414_/CLK _18955_/D vssd1 vssd1 vccd1 vccd1 _18955_/Q sky130_fd_sc_hd__dfxtp_1
X_14078_ _14078_/A _14078_/B vssd1 vssd1 vccd1 vccd1 _14078_/Y sky130_fd_sc_hd__nand2_1
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17906_ _12361_/A _17886_/X _12365_/X _12369_/X _17895_/X vssd1 vssd1 vccd1 vccd1
+ _19755_/D sky130_fd_sc_hd__o221a_1
X_13029_ _18321_/Q _13025_/C _13028_/Y vssd1 vssd1 vccd1 vccd1 _18321_/D sky130_fd_sc_hd__o21a_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18886_ _19703_/CLK _18886_/D vssd1 vssd1 vccd1 vccd1 _18886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17837_ _17837_/A vssd1 vssd1 vccd1 vccd1 _19719_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15084__A0 _18620_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17768_ _12193_/X _13423_/X _17625_/S vssd1 vssd1 vccd1 vccd1 _17768_/X sky130_fd_sc_hd__a21bo_1
XFILLER_54_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_75_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16719_ _19299_/Q _16718_/X _16719_/S vssd1 vssd1 vccd1 vccd1 _16720_/A sky130_fd_sc_hd__mux2_1
X_19507_ _19571_/CLK _19507_/D vssd1 vssd1 vccd1 vccd1 _19507_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09302__A2 _18533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17699_ _19676_/Q _17698_/X _17718_/S vssd1 vssd1 vccd1 vccd1 _17700_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19438_ _19699_/CLK _19438_/D vssd1 vssd1 vccd1 vccd1 _19438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19369_ _19550_/CLK _19369_/D vssd1 vssd1 vccd1 vccd1 _19369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16407__S _16413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14716__A _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09122_ _18554_/Q vssd1 vssd1 vccd1 vccd1 _11297_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15311__S _15311_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12070__A0 _12066_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13620__A _13620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17238__S _17241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16142__S _16150_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09955_ _09955_/A _18871_/Q vssd1 vssd1 vccd1 vccd1 _09955_/Y sky130_fd_sc_hd__nor2_1
XFILLER_132_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12125__A1 _19745_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15981__S _15983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10136__B1 _09621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ _09947_/A _09886_/B vssd1 vssd1 vccd1 vccd1 _09886_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10730_ _09408_/A _10716_/X _10721_/X _10729_/X _10846_/A vssd1 vssd1 vccd1 vccd1
+ _10730_/X sky130_fd_sc_hd__a221o_1
XANTENNA__15378__A1 _15191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14586__C1 _14585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10661_ _19691_/Q vssd1 vssd1 vccd1 vccd1 _10959_/A sky130_fd_sc_hd__buf_2
XFILLER_9_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14050__A1 _11899_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15221__S _15233_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12061__A0 _11135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12400_ _11200_/A _18519_/Q _12423_/S vssd1 vssd1 vccd1 vccd1 _12401_/A sky130_fd_sc_hd__mux2_8
X_13380_ _18294_/Q _13126_/X _13127_/X _18377_/Q vssd1 vssd1 vccd1 vccd1 _13380_/X
+ sky130_fd_sc_hd__a22o_1
X_10592_ _19638_/Q _19055_/Q _19092_/Q _18698_/Q _10511_/S _09515_/A vssd1 vssd1 vccd1
+ vccd1 _10593_/B sky130_fd_sc_hd__mux4_1
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10611__A1 _19187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14338__C1 _15116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12331_ _12285_/A _12309_/Y _12311_/B vssd1 vssd1 vccd1 vccd1 _12331_/X sky130_fd_sc_hd__o21a_1
XFILLER_127_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11688__C _11688_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15050_ _15048_/Y _15059_/B _14737_/A vssd1 vssd1 vccd1 vccd1 _15050_/Y sky130_fd_sc_hd__o21ai_1
X_12262_ _12262_/A _12262_/B vssd1 vssd1 vccd1 vccd1 _12265_/A sky130_fd_sc_hd__xnor2_4
XFILLER_119_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14001_ _13838_/A _13652_/X _13816_/A vssd1 vssd1 vccd1 vccd1 _14001_/Y sky130_fd_sc_hd__o21ai_1
X_11213_ _11551_/A _13526_/A _11299_/A vssd1 vssd1 vccd1 vccd1 _11213_/X sky130_fd_sc_hd__or3_1
X_12193_ _17143_/S vssd1 vssd1 vccd1 vccd1 _12193_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_123_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11144_ _12495_/C _09951_/A vssd1 vssd1 vccd1 vccd1 _11145_/A sky130_fd_sc_hd__or2b_1
XFILLER_122_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput74 _11926_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[10] sky130_fd_sc_hd__buf_2
Xoutput85 _12185_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[20] sky130_fd_sc_hd__buf_2
XFILLER_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput96 _12432_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[30] sky130_fd_sc_hd__buf_2
XANTENNA__15891__S _15891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18740_ _19616_/CLK _18740_/D vssd1 vssd1 vccd1 vccd1 _18740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11075_ _11075_/A _12468_/A vssd1 vssd1 vccd1 vccd1 _11254_/C sky130_fd_sc_hd__nor2_1
XFILLER_89_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15952_ _18207_/A _15952_/B vssd1 vssd1 vccd1 vccd1 _18977_/D sky130_fd_sc_hd__nor2_2
XANTENNA__10101__A_N _10098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10026_ _10020_/A _10023_/X _10025_/X _09988_/X vssd1 vssd1 vccd1 vccd1 _10026_/X
+ sky130_fd_sc_hd__o211a_1
X_14903_ _14903_/A _15000_/A vssd1 vssd1 vccd1 vccd1 _14925_/A sky130_fd_sc_hd__or2_1
X_18671_ _19326_/CLK _18671_/D vssd1 vssd1 vccd1 vccd1 _18671_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17391__B _17391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15883_ _14714_/X _18945_/Q _15891_/S vssd1 vssd1 vccd1 vccd1 _15884_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10773__S1 _10772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17622_ _17621_/A _17621_/C _14765_/A vssd1 vssd1 vccd1 vccd1 _17623_/B sky130_fd_sc_hd__o21ai_1
XFILLER_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14834_ _15077_/S vssd1 vssd1 vccd1 vccd1 _14880_/S sky130_fd_sc_hd__buf_2
XFILLER_56_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09190__A _09190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17553_ _19636_/Q _16768_/A _17557_/S vssd1 vssd1 vccd1 vccd1 _17554_/A sky130_fd_sc_hd__mux2_1
X_14765_ _14765_/A _18463_/Q _14765_/C vssd1 vssd1 vccd1 vccd1 _14786_/C sky130_fd_sc_hd__and3_1
XFILLER_147_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11977_ _11925_/A _11925_/B _11956_/A _11976_/Y vssd1 vssd1 vccd1 vccd1 _11978_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_16_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16504_ _16560_/A vssd1 vssd1 vccd1 vccd1 _16573_/S sky130_fd_sc_hd__buf_8
XFILLER_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13716_ _14332_/A vssd1 vssd1 vccd1 vccd1 _14285_/A sky130_fd_sc_hd__clkbuf_2
X_10928_ _10928_/A _10928_/B vssd1 vssd1 vccd1 vccd1 _10928_/X sky130_fd_sc_hd__or2_1
X_17484_ _17484_/A vssd1 vssd1 vccd1 vccd1 _19605_/D sky130_fd_sc_hd__clkbuf_1
X_14696_ _14696_/A vssd1 vssd1 vccd1 vccd1 _17890_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19223_ _19223_/CLK _19223_/D vssd1 vssd1 vccd1 vccd1 _19223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16435_ _16435_/A vssd1 vssd1 vccd1 vccd1 _19179_/D sky130_fd_sc_hd__clkbuf_1
X_13647_ _13665_/A _12401_/A _13659_/S vssd1 vssd1 vccd1 vccd1 _13647_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10859_ _09629_/A _10835_/Y _10858_/Y _10740_/X vssd1 vssd1 vccd1 vccd1 _10859_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19154_ _19702_/CLK _19154_/D vssd1 vssd1 vccd1 vccd1 _19154_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10289__S0 _09675_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _16366_/A vssd1 vssd1 vccd1 vccd1 _19149_/D sky130_fd_sc_hd__clkbuf_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _13578_/A _13584_/C _11599_/B _13545_/B vssd1 vssd1 vccd1 vccd1 _13579_/D
+ sky130_fd_sc_hd__or4bb_1
XANTENNA__11582__A1_N _18561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18105_ _18114_/A _18105_/B vssd1 vssd1 vccd1 vccd1 _18105_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15317_ _15317_/A vssd1 vssd1 vccd1 vccd1 _18710_/D sky130_fd_sc_hd__clkbuf_1
X_12529_ _12545_/A vssd1 vssd1 vccd1 vccd1 _12734_/A sky130_fd_sc_hd__buf_2
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19085_ _19633_/CLK _19085_/D vssd1 vssd1 vccd1 vccd1 _19085_/Q sky130_fd_sc_hd__dfxtp_1
X_16297_ _16297_/A vssd1 vssd1 vccd1 vccd1 _19119_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18036_ _18036_/A vssd1 vssd1 vccd1 vccd1 _18043_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_15248_ _17730_/A _13136_/X _11719_/B vssd1 vssd1 vccd1 vccd1 _15248_/X sky130_fd_sc_hd__a21o_1
XFILLER_114_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17058__S _17058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15179_ _18663_/Q _15178_/X _15185_/S vssd1 vssd1 vccd1 vccd1 _15180_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17294__A1 _16705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09740_ _10127_/A _09737_/X _09739_/X vssd1 vssd1 vccd1 vccd1 _09740_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_100_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18938_ _19556_/CLK _18938_/D vssd1 vssd1 vccd1 vccd1 _18938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
.ends

