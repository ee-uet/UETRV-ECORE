magic
tech sky130A
magscale 1 2
timestamp 1649143084
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 1104 2048 99898 97504
<< metal2 >>
rect 24950 99200 25006 100000
rect 74906 99200 74962 100000
rect 49974 0 50030 800
<< obsm2 >>
rect 1398 99144 24894 99657
rect 25062 99144 74850 99657
rect 75018 99144 99894 99657
rect 1398 856 99894 99144
rect 1398 303 49918 856
rect 50086 303 99894 856
<< metal3 >>
rect 99200 99560 100000 99680
rect 99200 99016 100000 99136
rect 99200 98472 100000 98592
rect 99200 97792 100000 97912
rect 99200 97248 100000 97368
rect 99200 96704 100000 96824
rect 99200 96160 100000 96280
rect 99200 95480 100000 95600
rect 99200 94936 100000 95056
rect 99200 94392 100000 94512
rect 99200 93712 100000 93832
rect 99200 93168 100000 93288
rect 99200 92624 100000 92744
rect 99200 92080 100000 92200
rect 99200 91400 100000 91520
rect 99200 90856 100000 90976
rect 99200 90312 100000 90432
rect 99200 89768 100000 89888
rect 99200 89088 100000 89208
rect 99200 88544 100000 88664
rect 99200 88000 100000 88120
rect 99200 87320 100000 87440
rect 99200 86776 100000 86896
rect 99200 86232 100000 86352
rect 99200 85688 100000 85808
rect 99200 85008 100000 85128
rect 99200 84464 100000 84584
rect 99200 83920 100000 84040
rect 99200 83376 100000 83496
rect 99200 82696 100000 82816
rect 99200 82152 100000 82272
rect 99200 81608 100000 81728
rect 99200 80928 100000 81048
rect 99200 80384 100000 80504
rect 99200 79840 100000 79960
rect 99200 79296 100000 79416
rect 99200 78616 100000 78736
rect 99200 78072 100000 78192
rect 99200 77528 100000 77648
rect 99200 76984 100000 77104
rect 99200 76304 100000 76424
rect 99200 75760 100000 75880
rect 99200 75216 100000 75336
rect 99200 74536 100000 74656
rect 99200 73992 100000 74112
rect 99200 73448 100000 73568
rect 99200 72904 100000 73024
rect 99200 72224 100000 72344
rect 99200 71680 100000 71800
rect 99200 71136 100000 71256
rect 99200 70592 100000 70712
rect 99200 69912 100000 70032
rect 99200 69368 100000 69488
rect 99200 68824 100000 68944
rect 99200 68144 100000 68264
rect 99200 67600 100000 67720
rect 99200 67056 100000 67176
rect 99200 66512 100000 66632
rect 99200 65832 100000 65952
rect 99200 65288 100000 65408
rect 99200 64744 100000 64864
rect 99200 64200 100000 64320
rect 99200 63520 100000 63640
rect 99200 62976 100000 63096
rect 99200 62432 100000 62552
rect 99200 61752 100000 61872
rect 99200 61208 100000 61328
rect 99200 60664 100000 60784
rect 99200 60120 100000 60240
rect 99200 59440 100000 59560
rect 99200 58896 100000 59016
rect 99200 58352 100000 58472
rect 99200 57808 100000 57928
rect 99200 57128 100000 57248
rect 99200 56584 100000 56704
rect 99200 56040 100000 56160
rect 99200 55360 100000 55480
rect 99200 54816 100000 54936
rect 99200 54272 100000 54392
rect 99200 53728 100000 53848
rect 99200 53048 100000 53168
rect 99200 52504 100000 52624
rect 99200 51960 100000 52080
rect 99200 51416 100000 51536
rect 99200 50736 100000 50856
rect 99200 50192 100000 50312
rect 0 49920 800 50040
rect 99200 49648 100000 49768
rect 99200 48968 100000 49088
rect 99200 48424 100000 48544
rect 99200 47880 100000 48000
rect 99200 47336 100000 47456
rect 99200 46656 100000 46776
rect 99200 46112 100000 46232
rect 99200 45568 100000 45688
rect 99200 45024 100000 45144
rect 99200 44344 100000 44464
rect 99200 43800 100000 43920
rect 99200 43256 100000 43376
rect 99200 42576 100000 42696
rect 99200 42032 100000 42152
rect 99200 41488 100000 41608
rect 99200 40944 100000 41064
rect 99200 40264 100000 40384
rect 99200 39720 100000 39840
rect 99200 39176 100000 39296
rect 99200 38632 100000 38752
rect 99200 37952 100000 38072
rect 99200 37408 100000 37528
rect 99200 36864 100000 36984
rect 99200 36184 100000 36304
rect 99200 35640 100000 35760
rect 99200 35096 100000 35216
rect 99200 34552 100000 34672
rect 99200 33872 100000 33992
rect 99200 33328 100000 33448
rect 99200 32784 100000 32904
rect 99200 32240 100000 32360
rect 99200 31560 100000 31680
rect 99200 31016 100000 31136
rect 99200 30472 100000 30592
rect 99200 29792 100000 29912
rect 99200 29248 100000 29368
rect 99200 28704 100000 28824
rect 99200 28160 100000 28280
rect 99200 27480 100000 27600
rect 99200 26936 100000 27056
rect 99200 26392 100000 26512
rect 99200 25848 100000 25968
rect 99200 25168 100000 25288
rect 99200 24624 100000 24744
rect 99200 24080 100000 24200
rect 99200 23400 100000 23520
rect 99200 22856 100000 22976
rect 99200 22312 100000 22432
rect 99200 21768 100000 21888
rect 99200 21088 100000 21208
rect 99200 20544 100000 20664
rect 99200 20000 100000 20120
rect 99200 19456 100000 19576
rect 99200 18776 100000 18896
rect 99200 18232 100000 18352
rect 99200 17688 100000 17808
rect 99200 17008 100000 17128
rect 99200 16464 100000 16584
rect 99200 15920 100000 16040
rect 99200 15376 100000 15496
rect 99200 14696 100000 14816
rect 99200 14152 100000 14272
rect 99200 13608 100000 13728
rect 99200 13064 100000 13184
rect 99200 12384 100000 12504
rect 99200 11840 100000 11960
rect 99200 11296 100000 11416
rect 99200 10616 100000 10736
rect 99200 10072 100000 10192
rect 99200 9528 100000 9648
rect 99200 8984 100000 9104
rect 99200 8304 100000 8424
rect 99200 7760 100000 7880
rect 99200 7216 100000 7336
rect 99200 6672 100000 6792
rect 99200 5992 100000 6112
rect 99200 5448 100000 5568
rect 99200 4904 100000 5024
rect 99200 4224 100000 4344
rect 99200 3680 100000 3800
rect 99200 3136 100000 3256
rect 99200 2592 100000 2712
rect 99200 1912 100000 2032
rect 99200 1368 100000 1488
rect 99200 824 100000 944
rect 99200 280 100000 400
<< obsm3 >>
rect 800 99480 99120 99653
rect 800 99216 99899 99480
rect 800 98936 99120 99216
rect 800 98672 99899 98936
rect 800 98392 99120 98672
rect 800 97992 99899 98392
rect 800 97712 99120 97992
rect 800 97448 99899 97712
rect 800 97168 99120 97448
rect 800 96904 99899 97168
rect 800 96624 99120 96904
rect 800 96360 99899 96624
rect 800 96080 99120 96360
rect 800 95680 99899 96080
rect 800 95400 99120 95680
rect 800 95136 99899 95400
rect 800 94856 99120 95136
rect 800 94592 99899 94856
rect 800 94312 99120 94592
rect 800 93912 99899 94312
rect 800 93632 99120 93912
rect 800 93368 99899 93632
rect 800 93088 99120 93368
rect 800 92824 99899 93088
rect 800 92544 99120 92824
rect 800 92280 99899 92544
rect 800 92000 99120 92280
rect 800 91600 99899 92000
rect 800 91320 99120 91600
rect 800 91056 99899 91320
rect 800 90776 99120 91056
rect 800 90512 99899 90776
rect 800 90232 99120 90512
rect 800 89968 99899 90232
rect 800 89688 99120 89968
rect 800 89288 99899 89688
rect 800 89008 99120 89288
rect 800 88744 99899 89008
rect 800 88464 99120 88744
rect 800 88200 99899 88464
rect 800 87920 99120 88200
rect 800 87520 99899 87920
rect 800 87240 99120 87520
rect 800 86976 99899 87240
rect 800 86696 99120 86976
rect 800 86432 99899 86696
rect 800 86152 99120 86432
rect 800 85888 99899 86152
rect 800 85608 99120 85888
rect 800 85208 99899 85608
rect 800 84928 99120 85208
rect 800 84664 99899 84928
rect 800 84384 99120 84664
rect 800 84120 99899 84384
rect 800 83840 99120 84120
rect 800 83576 99899 83840
rect 800 83296 99120 83576
rect 800 82896 99899 83296
rect 800 82616 99120 82896
rect 800 82352 99899 82616
rect 800 82072 99120 82352
rect 800 81808 99899 82072
rect 800 81528 99120 81808
rect 800 81128 99899 81528
rect 800 80848 99120 81128
rect 800 80584 99899 80848
rect 800 80304 99120 80584
rect 800 80040 99899 80304
rect 800 79760 99120 80040
rect 800 79496 99899 79760
rect 800 79216 99120 79496
rect 800 78816 99899 79216
rect 800 78536 99120 78816
rect 800 78272 99899 78536
rect 800 77992 99120 78272
rect 800 77728 99899 77992
rect 800 77448 99120 77728
rect 800 77184 99899 77448
rect 800 76904 99120 77184
rect 800 76504 99899 76904
rect 800 76224 99120 76504
rect 800 75960 99899 76224
rect 800 75680 99120 75960
rect 800 75416 99899 75680
rect 800 75136 99120 75416
rect 800 74736 99899 75136
rect 800 74456 99120 74736
rect 800 74192 99899 74456
rect 800 73912 99120 74192
rect 800 73648 99899 73912
rect 800 73368 99120 73648
rect 800 73104 99899 73368
rect 800 72824 99120 73104
rect 800 72424 99899 72824
rect 800 72144 99120 72424
rect 800 71880 99899 72144
rect 800 71600 99120 71880
rect 800 71336 99899 71600
rect 800 71056 99120 71336
rect 800 70792 99899 71056
rect 800 70512 99120 70792
rect 800 70112 99899 70512
rect 800 69832 99120 70112
rect 800 69568 99899 69832
rect 800 69288 99120 69568
rect 800 69024 99899 69288
rect 800 68744 99120 69024
rect 800 68344 99899 68744
rect 800 68064 99120 68344
rect 800 67800 99899 68064
rect 800 67520 99120 67800
rect 800 67256 99899 67520
rect 800 66976 99120 67256
rect 800 66712 99899 66976
rect 800 66432 99120 66712
rect 800 66032 99899 66432
rect 800 65752 99120 66032
rect 800 65488 99899 65752
rect 800 65208 99120 65488
rect 800 64944 99899 65208
rect 800 64664 99120 64944
rect 800 64400 99899 64664
rect 800 64120 99120 64400
rect 800 63720 99899 64120
rect 800 63440 99120 63720
rect 800 63176 99899 63440
rect 800 62896 99120 63176
rect 800 62632 99899 62896
rect 800 62352 99120 62632
rect 800 61952 99899 62352
rect 800 61672 99120 61952
rect 800 61408 99899 61672
rect 800 61128 99120 61408
rect 800 60864 99899 61128
rect 800 60584 99120 60864
rect 800 60320 99899 60584
rect 800 60040 99120 60320
rect 800 59640 99899 60040
rect 800 59360 99120 59640
rect 800 59096 99899 59360
rect 800 58816 99120 59096
rect 800 58552 99899 58816
rect 800 58272 99120 58552
rect 800 58008 99899 58272
rect 800 57728 99120 58008
rect 800 57328 99899 57728
rect 800 57048 99120 57328
rect 800 56784 99899 57048
rect 800 56504 99120 56784
rect 800 56240 99899 56504
rect 800 55960 99120 56240
rect 800 55560 99899 55960
rect 800 55280 99120 55560
rect 800 55016 99899 55280
rect 800 54736 99120 55016
rect 800 54472 99899 54736
rect 800 54192 99120 54472
rect 800 53928 99899 54192
rect 800 53648 99120 53928
rect 800 53248 99899 53648
rect 800 52968 99120 53248
rect 800 52704 99899 52968
rect 800 52424 99120 52704
rect 800 52160 99899 52424
rect 800 51880 99120 52160
rect 800 51616 99899 51880
rect 800 51336 99120 51616
rect 800 50936 99899 51336
rect 800 50656 99120 50936
rect 800 50392 99899 50656
rect 800 50120 99120 50392
rect 880 50112 99120 50120
rect 880 49848 99899 50112
rect 880 49840 99120 49848
rect 800 49568 99120 49840
rect 800 49168 99899 49568
rect 800 48888 99120 49168
rect 800 48624 99899 48888
rect 800 48344 99120 48624
rect 800 48080 99899 48344
rect 800 47800 99120 48080
rect 800 47536 99899 47800
rect 800 47256 99120 47536
rect 800 46856 99899 47256
rect 800 46576 99120 46856
rect 800 46312 99899 46576
rect 800 46032 99120 46312
rect 800 45768 99899 46032
rect 800 45488 99120 45768
rect 800 45224 99899 45488
rect 800 44944 99120 45224
rect 800 44544 99899 44944
rect 800 44264 99120 44544
rect 800 44000 99899 44264
rect 800 43720 99120 44000
rect 800 43456 99899 43720
rect 800 43176 99120 43456
rect 800 42776 99899 43176
rect 800 42496 99120 42776
rect 800 42232 99899 42496
rect 800 41952 99120 42232
rect 800 41688 99899 41952
rect 800 41408 99120 41688
rect 800 41144 99899 41408
rect 800 40864 99120 41144
rect 800 40464 99899 40864
rect 800 40184 99120 40464
rect 800 39920 99899 40184
rect 800 39640 99120 39920
rect 800 39376 99899 39640
rect 800 39096 99120 39376
rect 800 38832 99899 39096
rect 800 38552 99120 38832
rect 800 38152 99899 38552
rect 800 37872 99120 38152
rect 800 37608 99899 37872
rect 800 37328 99120 37608
rect 800 37064 99899 37328
rect 800 36784 99120 37064
rect 800 36384 99899 36784
rect 800 36104 99120 36384
rect 800 35840 99899 36104
rect 800 35560 99120 35840
rect 800 35296 99899 35560
rect 800 35016 99120 35296
rect 800 34752 99899 35016
rect 800 34472 99120 34752
rect 800 34072 99899 34472
rect 800 33792 99120 34072
rect 800 33528 99899 33792
rect 800 33248 99120 33528
rect 800 32984 99899 33248
rect 800 32704 99120 32984
rect 800 32440 99899 32704
rect 800 32160 99120 32440
rect 800 31760 99899 32160
rect 800 31480 99120 31760
rect 800 31216 99899 31480
rect 800 30936 99120 31216
rect 800 30672 99899 30936
rect 800 30392 99120 30672
rect 800 29992 99899 30392
rect 800 29712 99120 29992
rect 800 29448 99899 29712
rect 800 29168 99120 29448
rect 800 28904 99899 29168
rect 800 28624 99120 28904
rect 800 28360 99899 28624
rect 800 28080 99120 28360
rect 800 27680 99899 28080
rect 800 27400 99120 27680
rect 800 27136 99899 27400
rect 800 26856 99120 27136
rect 800 26592 99899 26856
rect 800 26312 99120 26592
rect 800 26048 99899 26312
rect 800 25768 99120 26048
rect 800 25368 99899 25768
rect 800 25088 99120 25368
rect 800 24824 99899 25088
rect 800 24544 99120 24824
rect 800 24280 99899 24544
rect 800 24000 99120 24280
rect 800 23600 99899 24000
rect 800 23320 99120 23600
rect 800 23056 99899 23320
rect 800 22776 99120 23056
rect 800 22512 99899 22776
rect 800 22232 99120 22512
rect 800 21968 99899 22232
rect 800 21688 99120 21968
rect 800 21288 99899 21688
rect 800 21008 99120 21288
rect 800 20744 99899 21008
rect 800 20464 99120 20744
rect 800 20200 99899 20464
rect 800 19920 99120 20200
rect 800 19656 99899 19920
rect 800 19376 99120 19656
rect 800 18976 99899 19376
rect 800 18696 99120 18976
rect 800 18432 99899 18696
rect 800 18152 99120 18432
rect 800 17888 99899 18152
rect 800 17608 99120 17888
rect 800 17208 99899 17608
rect 800 16928 99120 17208
rect 800 16664 99899 16928
rect 800 16384 99120 16664
rect 800 16120 99899 16384
rect 800 15840 99120 16120
rect 800 15576 99899 15840
rect 800 15296 99120 15576
rect 800 14896 99899 15296
rect 800 14616 99120 14896
rect 800 14352 99899 14616
rect 800 14072 99120 14352
rect 800 13808 99899 14072
rect 800 13528 99120 13808
rect 800 13264 99899 13528
rect 800 12984 99120 13264
rect 800 12584 99899 12984
rect 800 12304 99120 12584
rect 800 12040 99899 12304
rect 800 11760 99120 12040
rect 800 11496 99899 11760
rect 800 11216 99120 11496
rect 800 10816 99899 11216
rect 800 10536 99120 10816
rect 800 10272 99899 10536
rect 800 9992 99120 10272
rect 800 9728 99899 9992
rect 800 9448 99120 9728
rect 800 9184 99899 9448
rect 800 8904 99120 9184
rect 800 8504 99899 8904
rect 800 8224 99120 8504
rect 800 7960 99899 8224
rect 800 7680 99120 7960
rect 800 7416 99899 7680
rect 800 7136 99120 7416
rect 800 6872 99899 7136
rect 800 6592 99120 6872
rect 800 6192 99899 6592
rect 800 5912 99120 6192
rect 800 5648 99899 5912
rect 800 5368 99120 5648
rect 800 5104 99899 5368
rect 800 4824 99120 5104
rect 800 4424 99899 4824
rect 800 4144 99120 4424
rect 800 3880 99899 4144
rect 800 3600 99120 3880
rect 800 3336 99899 3600
rect 800 3056 99120 3336
rect 800 2792 99899 3056
rect 800 2512 99120 2792
rect 800 2112 99899 2512
rect 800 1832 99120 2112
rect 800 1568 99899 1832
rect 800 1288 99120 1568
rect 800 1024 99899 1288
rect 800 744 99120 1024
rect 800 480 99899 744
rect 800 307 99120 480
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< obsm4 >>
rect 3555 2347 4128 96661
rect 4608 2347 19488 96661
rect 19968 2347 34848 96661
rect 35328 2347 50208 96661
rect 50688 2347 65568 96661
rect 66048 2347 80928 96661
rect 81408 2347 96288 96661
rect 96768 2347 98197 96661
<< labels >>
rlabel metal2 s 24950 99200 25006 100000 6 clock
port 1 nsew signal input
rlabel metal3 s 99200 1912 100000 2032 6 io_dbus_addr[0]
port 2 nsew signal output
rlabel metal3 s 99200 22312 100000 22432 6 io_dbus_addr[10]
port 3 nsew signal output
rlabel metal3 s 99200 24080 100000 24200 6 io_dbus_addr[11]
port 4 nsew signal output
rlabel metal3 s 99200 25848 100000 25968 6 io_dbus_addr[12]
port 5 nsew signal output
rlabel metal3 s 99200 27480 100000 27600 6 io_dbus_addr[13]
port 6 nsew signal output
rlabel metal3 s 99200 29248 100000 29368 6 io_dbus_addr[14]
port 7 nsew signal output
rlabel metal3 s 99200 31016 100000 31136 6 io_dbus_addr[15]
port 8 nsew signal output
rlabel metal3 s 99200 32784 100000 32904 6 io_dbus_addr[16]
port 9 nsew signal output
rlabel metal3 s 99200 34552 100000 34672 6 io_dbus_addr[17]
port 10 nsew signal output
rlabel metal3 s 99200 36184 100000 36304 6 io_dbus_addr[18]
port 11 nsew signal output
rlabel metal3 s 99200 37952 100000 38072 6 io_dbus_addr[19]
port 12 nsew signal output
rlabel metal3 s 99200 4904 100000 5024 6 io_dbus_addr[1]
port 13 nsew signal output
rlabel metal3 s 99200 39720 100000 39840 6 io_dbus_addr[20]
port 14 nsew signal output
rlabel metal3 s 99200 41488 100000 41608 6 io_dbus_addr[21]
port 15 nsew signal output
rlabel metal3 s 99200 43256 100000 43376 6 io_dbus_addr[22]
port 16 nsew signal output
rlabel metal3 s 99200 45024 100000 45144 6 io_dbus_addr[23]
port 17 nsew signal output
rlabel metal3 s 99200 46656 100000 46776 6 io_dbus_addr[24]
port 18 nsew signal output
rlabel metal3 s 99200 48424 100000 48544 6 io_dbus_addr[25]
port 19 nsew signal output
rlabel metal3 s 99200 50192 100000 50312 6 io_dbus_addr[26]
port 20 nsew signal output
rlabel metal3 s 99200 51960 100000 52080 6 io_dbus_addr[27]
port 21 nsew signal output
rlabel metal3 s 99200 53728 100000 53848 6 io_dbus_addr[28]
port 22 nsew signal output
rlabel metal3 s 99200 55360 100000 55480 6 io_dbus_addr[29]
port 23 nsew signal output
rlabel metal3 s 99200 7760 100000 7880 6 io_dbus_addr[2]
port 24 nsew signal output
rlabel metal3 s 99200 57128 100000 57248 6 io_dbus_addr[30]
port 25 nsew signal output
rlabel metal3 s 99200 58896 100000 59016 6 io_dbus_addr[31]
port 26 nsew signal output
rlabel metal3 s 99200 10072 100000 10192 6 io_dbus_addr[3]
port 27 nsew signal output
rlabel metal3 s 99200 11840 100000 11960 6 io_dbus_addr[4]
port 28 nsew signal output
rlabel metal3 s 99200 13608 100000 13728 6 io_dbus_addr[5]
port 29 nsew signal output
rlabel metal3 s 99200 15376 100000 15496 6 io_dbus_addr[6]
port 30 nsew signal output
rlabel metal3 s 99200 17008 100000 17128 6 io_dbus_addr[7]
port 31 nsew signal output
rlabel metal3 s 99200 18776 100000 18896 6 io_dbus_addr[8]
port 32 nsew signal output
rlabel metal3 s 99200 20544 100000 20664 6 io_dbus_addr[9]
port 33 nsew signal output
rlabel metal3 s 99200 2592 100000 2712 6 io_dbus_ld_type[0]
port 34 nsew signal output
rlabel metal3 s 99200 5448 100000 5568 6 io_dbus_ld_type[1]
port 35 nsew signal output
rlabel metal3 s 99200 8304 100000 8424 6 io_dbus_ld_type[2]
port 36 nsew signal output
rlabel metal3 s 99200 280 100000 400 6 io_dbus_rd_en
port 37 nsew signal output
rlabel metal3 s 99200 3136 100000 3256 6 io_dbus_rdata[0]
port 38 nsew signal input
rlabel metal3 s 99200 22856 100000 22976 6 io_dbus_rdata[10]
port 39 nsew signal input
rlabel metal3 s 99200 24624 100000 24744 6 io_dbus_rdata[11]
port 40 nsew signal input
rlabel metal3 s 99200 26392 100000 26512 6 io_dbus_rdata[12]
port 41 nsew signal input
rlabel metal3 s 99200 28160 100000 28280 6 io_dbus_rdata[13]
port 42 nsew signal input
rlabel metal3 s 99200 29792 100000 29912 6 io_dbus_rdata[14]
port 43 nsew signal input
rlabel metal3 s 99200 31560 100000 31680 6 io_dbus_rdata[15]
port 44 nsew signal input
rlabel metal3 s 99200 33328 100000 33448 6 io_dbus_rdata[16]
port 45 nsew signal input
rlabel metal3 s 99200 35096 100000 35216 6 io_dbus_rdata[17]
port 46 nsew signal input
rlabel metal3 s 99200 36864 100000 36984 6 io_dbus_rdata[18]
port 47 nsew signal input
rlabel metal3 s 99200 38632 100000 38752 6 io_dbus_rdata[19]
port 48 nsew signal input
rlabel metal3 s 99200 5992 100000 6112 6 io_dbus_rdata[1]
port 49 nsew signal input
rlabel metal3 s 99200 40264 100000 40384 6 io_dbus_rdata[20]
port 50 nsew signal input
rlabel metal3 s 99200 42032 100000 42152 6 io_dbus_rdata[21]
port 51 nsew signal input
rlabel metal3 s 99200 43800 100000 43920 6 io_dbus_rdata[22]
port 52 nsew signal input
rlabel metal3 s 99200 45568 100000 45688 6 io_dbus_rdata[23]
port 53 nsew signal input
rlabel metal3 s 99200 47336 100000 47456 6 io_dbus_rdata[24]
port 54 nsew signal input
rlabel metal3 s 99200 48968 100000 49088 6 io_dbus_rdata[25]
port 55 nsew signal input
rlabel metal3 s 99200 50736 100000 50856 6 io_dbus_rdata[26]
port 56 nsew signal input
rlabel metal3 s 99200 52504 100000 52624 6 io_dbus_rdata[27]
port 57 nsew signal input
rlabel metal3 s 99200 54272 100000 54392 6 io_dbus_rdata[28]
port 58 nsew signal input
rlabel metal3 s 99200 56040 100000 56160 6 io_dbus_rdata[29]
port 59 nsew signal input
rlabel metal3 s 99200 8984 100000 9104 6 io_dbus_rdata[2]
port 60 nsew signal input
rlabel metal3 s 99200 57808 100000 57928 6 io_dbus_rdata[30]
port 61 nsew signal input
rlabel metal3 s 99200 59440 100000 59560 6 io_dbus_rdata[31]
port 62 nsew signal input
rlabel metal3 s 99200 10616 100000 10736 6 io_dbus_rdata[3]
port 63 nsew signal input
rlabel metal3 s 99200 12384 100000 12504 6 io_dbus_rdata[4]
port 64 nsew signal input
rlabel metal3 s 99200 14152 100000 14272 6 io_dbus_rdata[5]
port 65 nsew signal input
rlabel metal3 s 99200 15920 100000 16040 6 io_dbus_rdata[6]
port 66 nsew signal input
rlabel metal3 s 99200 17688 100000 17808 6 io_dbus_rdata[7]
port 67 nsew signal input
rlabel metal3 s 99200 19456 100000 19576 6 io_dbus_rdata[8]
port 68 nsew signal input
rlabel metal3 s 99200 21088 100000 21208 6 io_dbus_rdata[9]
port 69 nsew signal input
rlabel metal3 s 99200 3680 100000 3800 6 io_dbus_st_type[0]
port 70 nsew signal output
rlabel metal3 s 99200 6672 100000 6792 6 io_dbus_st_type[1]
port 71 nsew signal output
rlabel metal3 s 99200 824 100000 944 6 io_dbus_valid
port 72 nsew signal input
rlabel metal3 s 99200 4224 100000 4344 6 io_dbus_wdata[0]
port 73 nsew signal output
rlabel metal3 s 99200 23400 100000 23520 6 io_dbus_wdata[10]
port 74 nsew signal output
rlabel metal3 s 99200 25168 100000 25288 6 io_dbus_wdata[11]
port 75 nsew signal output
rlabel metal3 s 99200 26936 100000 27056 6 io_dbus_wdata[12]
port 76 nsew signal output
rlabel metal3 s 99200 28704 100000 28824 6 io_dbus_wdata[13]
port 77 nsew signal output
rlabel metal3 s 99200 30472 100000 30592 6 io_dbus_wdata[14]
port 78 nsew signal output
rlabel metal3 s 99200 32240 100000 32360 6 io_dbus_wdata[15]
port 79 nsew signal output
rlabel metal3 s 99200 33872 100000 33992 6 io_dbus_wdata[16]
port 80 nsew signal output
rlabel metal3 s 99200 35640 100000 35760 6 io_dbus_wdata[17]
port 81 nsew signal output
rlabel metal3 s 99200 37408 100000 37528 6 io_dbus_wdata[18]
port 82 nsew signal output
rlabel metal3 s 99200 39176 100000 39296 6 io_dbus_wdata[19]
port 83 nsew signal output
rlabel metal3 s 99200 7216 100000 7336 6 io_dbus_wdata[1]
port 84 nsew signal output
rlabel metal3 s 99200 40944 100000 41064 6 io_dbus_wdata[20]
port 85 nsew signal output
rlabel metal3 s 99200 42576 100000 42696 6 io_dbus_wdata[21]
port 86 nsew signal output
rlabel metal3 s 99200 44344 100000 44464 6 io_dbus_wdata[22]
port 87 nsew signal output
rlabel metal3 s 99200 46112 100000 46232 6 io_dbus_wdata[23]
port 88 nsew signal output
rlabel metal3 s 99200 47880 100000 48000 6 io_dbus_wdata[24]
port 89 nsew signal output
rlabel metal3 s 99200 49648 100000 49768 6 io_dbus_wdata[25]
port 90 nsew signal output
rlabel metal3 s 99200 51416 100000 51536 6 io_dbus_wdata[26]
port 91 nsew signal output
rlabel metal3 s 99200 53048 100000 53168 6 io_dbus_wdata[27]
port 92 nsew signal output
rlabel metal3 s 99200 54816 100000 54936 6 io_dbus_wdata[28]
port 93 nsew signal output
rlabel metal3 s 99200 56584 100000 56704 6 io_dbus_wdata[29]
port 94 nsew signal output
rlabel metal3 s 99200 9528 100000 9648 6 io_dbus_wdata[2]
port 95 nsew signal output
rlabel metal3 s 99200 58352 100000 58472 6 io_dbus_wdata[30]
port 96 nsew signal output
rlabel metal3 s 99200 60120 100000 60240 6 io_dbus_wdata[31]
port 97 nsew signal output
rlabel metal3 s 99200 11296 100000 11416 6 io_dbus_wdata[3]
port 98 nsew signal output
rlabel metal3 s 99200 13064 100000 13184 6 io_dbus_wdata[4]
port 99 nsew signal output
rlabel metal3 s 99200 14696 100000 14816 6 io_dbus_wdata[5]
port 100 nsew signal output
rlabel metal3 s 99200 16464 100000 16584 6 io_dbus_wdata[6]
port 101 nsew signal output
rlabel metal3 s 99200 18232 100000 18352 6 io_dbus_wdata[7]
port 102 nsew signal output
rlabel metal3 s 99200 20000 100000 20120 6 io_dbus_wdata[8]
port 103 nsew signal output
rlabel metal3 s 99200 21768 100000 21888 6 io_dbus_wdata[9]
port 104 nsew signal output
rlabel metal3 s 99200 1368 100000 1488 6 io_dbus_wr_en
port 105 nsew signal output
rlabel metal3 s 99200 61208 100000 61328 6 io_ibus_addr[0]
port 106 nsew signal output
rlabel metal3 s 99200 72904 100000 73024 6 io_ibus_addr[10]
port 107 nsew signal output
rlabel metal3 s 99200 73992 100000 74112 6 io_ibus_addr[11]
port 108 nsew signal output
rlabel metal3 s 99200 75216 100000 75336 6 io_ibus_addr[12]
port 109 nsew signal output
rlabel metal3 s 99200 76304 100000 76424 6 io_ibus_addr[13]
port 110 nsew signal output
rlabel metal3 s 99200 77528 100000 77648 6 io_ibus_addr[14]
port 111 nsew signal output
rlabel metal3 s 99200 78616 100000 78736 6 io_ibus_addr[15]
port 112 nsew signal output
rlabel metal3 s 99200 79840 100000 79960 6 io_ibus_addr[16]
port 113 nsew signal output
rlabel metal3 s 99200 80928 100000 81048 6 io_ibus_addr[17]
port 114 nsew signal output
rlabel metal3 s 99200 82152 100000 82272 6 io_ibus_addr[18]
port 115 nsew signal output
rlabel metal3 s 99200 83376 100000 83496 6 io_ibus_addr[19]
port 116 nsew signal output
rlabel metal3 s 99200 62432 100000 62552 6 io_ibus_addr[1]
port 117 nsew signal output
rlabel metal3 s 99200 84464 100000 84584 6 io_ibus_addr[20]
port 118 nsew signal output
rlabel metal3 s 99200 85688 100000 85808 6 io_ibus_addr[21]
port 119 nsew signal output
rlabel metal3 s 99200 86776 100000 86896 6 io_ibus_addr[22]
port 120 nsew signal output
rlabel metal3 s 99200 88000 100000 88120 6 io_ibus_addr[23]
port 121 nsew signal output
rlabel metal3 s 99200 89088 100000 89208 6 io_ibus_addr[24]
port 122 nsew signal output
rlabel metal3 s 99200 90312 100000 90432 6 io_ibus_addr[25]
port 123 nsew signal output
rlabel metal3 s 99200 91400 100000 91520 6 io_ibus_addr[26]
port 124 nsew signal output
rlabel metal3 s 99200 92624 100000 92744 6 io_ibus_addr[27]
port 125 nsew signal output
rlabel metal3 s 99200 93712 100000 93832 6 io_ibus_addr[28]
port 126 nsew signal output
rlabel metal3 s 99200 94936 100000 95056 6 io_ibus_addr[29]
port 127 nsew signal output
rlabel metal3 s 99200 63520 100000 63640 6 io_ibus_addr[2]
port 128 nsew signal output
rlabel metal3 s 99200 96160 100000 96280 6 io_ibus_addr[30]
port 129 nsew signal output
rlabel metal3 s 99200 97248 100000 97368 6 io_ibus_addr[31]
port 130 nsew signal output
rlabel metal3 s 99200 64744 100000 64864 6 io_ibus_addr[3]
port 131 nsew signal output
rlabel metal3 s 99200 65832 100000 65952 6 io_ibus_addr[4]
port 132 nsew signal output
rlabel metal3 s 99200 67056 100000 67176 6 io_ibus_addr[5]
port 133 nsew signal output
rlabel metal3 s 99200 68144 100000 68264 6 io_ibus_addr[6]
port 134 nsew signal output
rlabel metal3 s 99200 69368 100000 69488 6 io_ibus_addr[7]
port 135 nsew signal output
rlabel metal3 s 99200 70592 100000 70712 6 io_ibus_addr[8]
port 136 nsew signal output
rlabel metal3 s 99200 71680 100000 71800 6 io_ibus_addr[9]
port 137 nsew signal output
rlabel metal3 s 99200 61752 100000 61872 6 io_ibus_inst[0]
port 138 nsew signal input
rlabel metal3 s 99200 73448 100000 73568 6 io_ibus_inst[10]
port 139 nsew signal input
rlabel metal3 s 99200 74536 100000 74656 6 io_ibus_inst[11]
port 140 nsew signal input
rlabel metal3 s 99200 75760 100000 75880 6 io_ibus_inst[12]
port 141 nsew signal input
rlabel metal3 s 99200 76984 100000 77104 6 io_ibus_inst[13]
port 142 nsew signal input
rlabel metal3 s 99200 78072 100000 78192 6 io_ibus_inst[14]
port 143 nsew signal input
rlabel metal3 s 99200 79296 100000 79416 6 io_ibus_inst[15]
port 144 nsew signal input
rlabel metal3 s 99200 80384 100000 80504 6 io_ibus_inst[16]
port 145 nsew signal input
rlabel metal3 s 99200 81608 100000 81728 6 io_ibus_inst[17]
port 146 nsew signal input
rlabel metal3 s 99200 82696 100000 82816 6 io_ibus_inst[18]
port 147 nsew signal input
rlabel metal3 s 99200 83920 100000 84040 6 io_ibus_inst[19]
port 148 nsew signal input
rlabel metal3 s 99200 62976 100000 63096 6 io_ibus_inst[1]
port 149 nsew signal input
rlabel metal3 s 99200 85008 100000 85128 6 io_ibus_inst[20]
port 150 nsew signal input
rlabel metal3 s 99200 86232 100000 86352 6 io_ibus_inst[21]
port 151 nsew signal input
rlabel metal3 s 99200 87320 100000 87440 6 io_ibus_inst[22]
port 152 nsew signal input
rlabel metal3 s 99200 88544 100000 88664 6 io_ibus_inst[23]
port 153 nsew signal input
rlabel metal3 s 99200 89768 100000 89888 6 io_ibus_inst[24]
port 154 nsew signal input
rlabel metal3 s 99200 90856 100000 90976 6 io_ibus_inst[25]
port 155 nsew signal input
rlabel metal3 s 99200 92080 100000 92200 6 io_ibus_inst[26]
port 156 nsew signal input
rlabel metal3 s 99200 93168 100000 93288 6 io_ibus_inst[27]
port 157 nsew signal input
rlabel metal3 s 99200 94392 100000 94512 6 io_ibus_inst[28]
port 158 nsew signal input
rlabel metal3 s 99200 95480 100000 95600 6 io_ibus_inst[29]
port 159 nsew signal input
rlabel metal3 s 99200 64200 100000 64320 6 io_ibus_inst[2]
port 160 nsew signal input
rlabel metal3 s 99200 96704 100000 96824 6 io_ibus_inst[30]
port 161 nsew signal input
rlabel metal3 s 99200 97792 100000 97912 6 io_ibus_inst[31]
port 162 nsew signal input
rlabel metal3 s 99200 65288 100000 65408 6 io_ibus_inst[3]
port 163 nsew signal input
rlabel metal3 s 99200 66512 100000 66632 6 io_ibus_inst[4]
port 164 nsew signal input
rlabel metal3 s 99200 67600 100000 67720 6 io_ibus_inst[5]
port 165 nsew signal input
rlabel metal3 s 99200 68824 100000 68944 6 io_ibus_inst[6]
port 166 nsew signal input
rlabel metal3 s 99200 69912 100000 70032 6 io_ibus_inst[7]
port 167 nsew signal input
rlabel metal3 s 99200 71136 100000 71256 6 io_ibus_inst[8]
port 168 nsew signal input
rlabel metal3 s 99200 72224 100000 72344 6 io_ibus_inst[9]
port 169 nsew signal input
rlabel metal3 s 99200 60664 100000 60784 6 io_ibus_valid
port 170 nsew signal input
rlabel metal3 s 99200 99560 100000 99680 6 io_irq_m1_irq
port 171 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 io_irq_m2_irq
port 172 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 io_irq_m3_irq
port 173 nsew signal input
rlabel metal3 s 99200 98472 100000 98592 6 io_irq_spi_irq
port 174 nsew signal input
rlabel metal3 s 99200 99016 100000 99136 6 io_irq_uart_irq
port 175 nsew signal input
rlabel metal2 s 74906 99200 74962 100000 6 reset
port 176 nsew signal input
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 177 nsew power input
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 177 nsew power input
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 177 nsew power input
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 177 nsew power input
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 178 nsew ground input
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 178 nsew ground input
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 178 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 35440734
string GDS_FILE /home/ali112000/Desktop/mpw/UETRV-ECORE/openlane/Core/runs/Core/results/finishing/Core.magic.gds
string GDS_START 1356826
<< end >>

