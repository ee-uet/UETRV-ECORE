magic
tech sky130A
magscale 1 2
timestamp 1647772013
<< obsli1 >>
rect 1104 2159 138828 137649
<< obsm1 >>
rect 1026 2128 139366 137828
<< metal2 >>
rect 662 139200 718 140000
rect 1950 139200 2006 140000
rect 3238 139200 3294 140000
rect 4526 139200 4582 140000
rect 5814 139200 5870 140000
rect 7102 139200 7158 140000
rect 8390 139200 8446 140000
rect 9678 139200 9734 140000
rect 10966 139200 11022 140000
rect 12254 139200 12310 140000
rect 13542 139200 13598 140000
rect 14922 139200 14978 140000
rect 16210 139200 16266 140000
rect 17498 139200 17554 140000
rect 18786 139200 18842 140000
rect 20074 139200 20130 140000
rect 21362 139200 21418 140000
rect 22650 139200 22706 140000
rect 23938 139200 23994 140000
rect 25226 139200 25282 140000
rect 26514 139200 26570 140000
rect 27802 139200 27858 140000
rect 29182 139200 29238 140000
rect 30470 139200 30526 140000
rect 31758 139200 31814 140000
rect 33046 139200 33102 140000
rect 34334 139200 34390 140000
rect 35622 139200 35678 140000
rect 36910 139200 36966 140000
rect 38198 139200 38254 140000
rect 39486 139200 39542 140000
rect 40774 139200 40830 140000
rect 42062 139200 42118 140000
rect 43442 139200 43498 140000
rect 44730 139200 44786 140000
rect 46018 139200 46074 140000
rect 47306 139200 47362 140000
rect 48594 139200 48650 140000
rect 49882 139200 49938 140000
rect 51170 139200 51226 140000
rect 52458 139200 52514 140000
rect 53746 139200 53802 140000
rect 55034 139200 55090 140000
rect 56322 139200 56378 140000
rect 57702 139200 57758 140000
rect 58990 139200 59046 140000
rect 60278 139200 60334 140000
rect 61566 139200 61622 140000
rect 62854 139200 62910 140000
rect 64142 139200 64198 140000
rect 65430 139200 65486 140000
rect 66718 139200 66774 140000
rect 68006 139200 68062 140000
rect 69294 139200 69350 140000
rect 70674 139200 70730 140000
rect 71962 139200 72018 140000
rect 73250 139200 73306 140000
rect 74538 139200 74594 140000
rect 75826 139200 75882 140000
rect 77114 139200 77170 140000
rect 78402 139200 78458 140000
rect 79690 139200 79746 140000
rect 80978 139200 81034 140000
rect 82266 139200 82322 140000
rect 83554 139200 83610 140000
rect 84934 139200 84990 140000
rect 86222 139200 86278 140000
rect 87510 139200 87566 140000
rect 88798 139200 88854 140000
rect 90086 139200 90142 140000
rect 91374 139200 91430 140000
rect 92662 139200 92718 140000
rect 93950 139200 94006 140000
rect 95238 139200 95294 140000
rect 96526 139200 96582 140000
rect 97814 139200 97870 140000
rect 99194 139200 99250 140000
rect 100482 139200 100538 140000
rect 101770 139200 101826 140000
rect 103058 139200 103114 140000
rect 104346 139200 104402 140000
rect 105634 139200 105690 140000
rect 106922 139200 106978 140000
rect 108210 139200 108266 140000
rect 109498 139200 109554 140000
rect 110786 139200 110842 140000
rect 112074 139200 112130 140000
rect 113454 139200 113510 140000
rect 114742 139200 114798 140000
rect 116030 139200 116086 140000
rect 117318 139200 117374 140000
rect 118606 139200 118662 140000
rect 119894 139200 119950 140000
rect 121182 139200 121238 140000
rect 122470 139200 122526 140000
rect 123758 139200 123814 140000
rect 125046 139200 125102 140000
rect 126334 139200 126390 140000
rect 127714 139200 127770 140000
rect 129002 139200 129058 140000
rect 130290 139200 130346 140000
rect 131578 139200 131634 140000
rect 132866 139200 132922 140000
rect 134154 139200 134210 140000
rect 135442 139200 135498 140000
rect 136730 139200 136786 140000
rect 138018 139200 138074 140000
rect 139306 139200 139362 140000
rect 3514 0 3570 800
rect 10506 0 10562 800
rect 17498 0 17554 800
rect 24490 0 24546 800
rect 31482 0 31538 800
rect 38474 0 38530 800
rect 45466 0 45522 800
rect 52458 0 52514 800
rect 59450 0 59506 800
rect 66442 0 66498 800
rect 73526 0 73582 800
rect 80518 0 80574 800
rect 87510 0 87566 800
rect 94502 0 94558 800
rect 101494 0 101550 800
rect 108486 0 108542 800
rect 115478 0 115534 800
rect 122470 0 122526 800
rect 129462 0 129518 800
rect 136454 0 136510 800
<< obsm2 >>
rect 774 139144 1894 139505
rect 2062 139144 3182 139505
rect 3350 139144 4470 139505
rect 4638 139144 5758 139505
rect 5926 139144 7046 139505
rect 7214 139144 8334 139505
rect 8502 139144 9622 139505
rect 9790 139144 10910 139505
rect 11078 139144 12198 139505
rect 12366 139144 13486 139505
rect 13654 139144 14866 139505
rect 15034 139144 16154 139505
rect 16322 139144 17442 139505
rect 17610 139144 18730 139505
rect 18898 139144 20018 139505
rect 20186 139144 21306 139505
rect 21474 139144 22594 139505
rect 22762 139144 23882 139505
rect 24050 139144 25170 139505
rect 25338 139144 26458 139505
rect 26626 139144 27746 139505
rect 27914 139144 29126 139505
rect 29294 139144 30414 139505
rect 30582 139144 31702 139505
rect 31870 139144 32990 139505
rect 33158 139144 34278 139505
rect 34446 139144 35566 139505
rect 35734 139144 36854 139505
rect 37022 139144 38142 139505
rect 38310 139144 39430 139505
rect 39598 139144 40718 139505
rect 40886 139144 42006 139505
rect 42174 139144 43386 139505
rect 43554 139144 44674 139505
rect 44842 139144 45962 139505
rect 46130 139144 47250 139505
rect 47418 139144 48538 139505
rect 48706 139144 49826 139505
rect 49994 139144 51114 139505
rect 51282 139144 52402 139505
rect 52570 139144 53690 139505
rect 53858 139144 54978 139505
rect 55146 139144 56266 139505
rect 56434 139144 57646 139505
rect 57814 139144 58934 139505
rect 59102 139144 60222 139505
rect 60390 139144 61510 139505
rect 61678 139144 62798 139505
rect 62966 139144 64086 139505
rect 64254 139144 65374 139505
rect 65542 139144 66662 139505
rect 66830 139144 67950 139505
rect 68118 139144 69238 139505
rect 69406 139144 70618 139505
rect 70786 139144 71906 139505
rect 72074 139144 73194 139505
rect 73362 139144 74482 139505
rect 74650 139144 75770 139505
rect 75938 139144 77058 139505
rect 77226 139144 78346 139505
rect 78514 139144 79634 139505
rect 79802 139144 80922 139505
rect 81090 139144 82210 139505
rect 82378 139144 83498 139505
rect 83666 139144 84878 139505
rect 85046 139144 86166 139505
rect 86334 139144 87454 139505
rect 87622 139144 88742 139505
rect 88910 139144 90030 139505
rect 90198 139144 91318 139505
rect 91486 139144 92606 139505
rect 92774 139144 93894 139505
rect 94062 139144 95182 139505
rect 95350 139144 96470 139505
rect 96638 139144 97758 139505
rect 97926 139144 99138 139505
rect 99306 139144 100426 139505
rect 100594 139144 101714 139505
rect 101882 139144 103002 139505
rect 103170 139144 104290 139505
rect 104458 139144 105578 139505
rect 105746 139144 106866 139505
rect 107034 139144 108154 139505
rect 108322 139144 109442 139505
rect 109610 139144 110730 139505
rect 110898 139144 112018 139505
rect 112186 139144 113398 139505
rect 113566 139144 114686 139505
rect 114854 139144 115974 139505
rect 116142 139144 117262 139505
rect 117430 139144 118550 139505
rect 118718 139144 119838 139505
rect 120006 139144 121126 139505
rect 121294 139144 122414 139505
rect 122582 139144 123702 139505
rect 123870 139144 124990 139505
rect 125158 139144 126278 139505
rect 126446 139144 127658 139505
rect 127826 139144 128946 139505
rect 129114 139144 130234 139505
rect 130402 139144 131522 139505
rect 131690 139144 132810 139505
rect 132978 139144 134098 139505
rect 134266 139144 135386 139505
rect 135554 139144 136674 139505
rect 136842 139144 137962 139505
rect 138130 139144 139250 139505
rect 718 856 139360 139144
rect 718 303 3458 856
rect 3626 303 10450 856
rect 10618 303 17442 856
rect 17610 303 24434 856
rect 24602 303 31426 856
rect 31594 303 38418 856
rect 38586 303 45410 856
rect 45578 303 52402 856
rect 52570 303 59394 856
rect 59562 303 66386 856
rect 66554 303 73470 856
rect 73638 303 80462 856
rect 80630 303 87454 856
rect 87622 303 94446 856
rect 94614 303 101438 856
rect 101606 303 108430 856
rect 108598 303 115422 856
rect 115590 303 122414 856
rect 122582 303 129406 856
rect 129574 303 136398 856
rect 136566 303 139360 856
<< metal3 >>
rect 0 139408 800 139528
rect 139200 139136 140000 139256
rect 0 138592 800 138712
rect 0 137912 800 138032
rect 139200 137912 140000 138032
rect 0 137096 800 137216
rect 139200 136552 140000 136672
rect 0 136280 800 136400
rect 0 135600 800 135720
rect 139200 135328 140000 135448
rect 0 134784 800 134904
rect 0 133968 800 134088
rect 139200 134104 140000 134224
rect 0 133288 800 133408
rect 139200 132744 140000 132864
rect 0 132472 800 132592
rect 0 131656 800 131776
rect 139200 131520 140000 131640
rect 0 130976 800 131096
rect 0 130160 800 130280
rect 139200 130296 140000 130416
rect 0 129344 800 129464
rect 139200 128936 140000 129056
rect 0 128664 800 128784
rect 0 127848 800 127968
rect 139200 127712 140000 127832
rect 0 127032 800 127152
rect 0 126352 800 126472
rect 139200 126488 140000 126608
rect 0 125536 800 125656
rect 139200 125128 140000 125248
rect 0 124720 800 124840
rect 0 124040 800 124160
rect 139200 123904 140000 124024
rect 0 123224 800 123344
rect 139200 122680 140000 122800
rect 0 122408 800 122528
rect 0 121728 800 121848
rect 139200 121320 140000 121440
rect 0 120912 800 121032
rect 0 120232 800 120352
rect 139200 120096 140000 120216
rect 0 119416 800 119536
rect 0 118600 800 118720
rect 139200 118736 140000 118856
rect 0 117920 800 118040
rect 139200 117512 140000 117632
rect 0 117104 800 117224
rect 0 116288 800 116408
rect 139200 116288 140000 116408
rect 0 115608 800 115728
rect 0 114792 800 114912
rect 139200 114928 140000 115048
rect 0 113976 800 114096
rect 139200 113704 140000 113824
rect 0 113296 800 113416
rect 0 112480 800 112600
rect 139200 112480 140000 112600
rect 0 111664 800 111784
rect 0 110984 800 111104
rect 139200 111120 140000 111240
rect 0 110168 800 110288
rect 139200 109896 140000 110016
rect 0 109352 800 109472
rect 0 108672 800 108792
rect 139200 108672 140000 108792
rect 0 107856 800 107976
rect 139200 107312 140000 107432
rect 0 107040 800 107160
rect 0 106360 800 106480
rect 139200 106088 140000 106208
rect 0 105544 800 105664
rect 0 104728 800 104848
rect 139200 104864 140000 104984
rect 0 104048 800 104168
rect 139200 103504 140000 103624
rect 0 103232 800 103352
rect 0 102416 800 102536
rect 139200 102280 140000 102400
rect 0 101736 800 101856
rect 0 100920 800 101040
rect 139200 101056 140000 101176
rect 0 100240 800 100360
rect 139200 99696 140000 99816
rect 0 99424 800 99544
rect 0 98608 800 98728
rect 139200 98472 140000 98592
rect 0 97928 800 98048
rect 0 97112 800 97232
rect 139200 97112 140000 97232
rect 0 96296 800 96416
rect 139200 95888 140000 96008
rect 0 95616 800 95736
rect 0 94800 800 94920
rect 139200 94664 140000 94784
rect 0 93984 800 94104
rect 0 93304 800 93424
rect 139200 93304 140000 93424
rect 0 92488 800 92608
rect 139200 92080 140000 92200
rect 0 91672 800 91792
rect 0 90992 800 91112
rect 139200 90856 140000 90976
rect 0 90176 800 90296
rect 0 89360 800 89480
rect 139200 89496 140000 89616
rect 0 88680 800 88800
rect 139200 88272 140000 88392
rect 0 87864 800 87984
rect 0 87048 800 87168
rect 139200 87048 140000 87168
rect 0 86368 800 86488
rect 0 85552 800 85672
rect 139200 85688 140000 85808
rect 0 84736 800 84856
rect 139200 84464 140000 84584
rect 0 84056 800 84176
rect 0 83240 800 83360
rect 139200 83240 140000 83360
rect 0 82424 800 82544
rect 0 81744 800 81864
rect 139200 81880 140000 82000
rect 0 80928 800 81048
rect 139200 80656 140000 80776
rect 0 80248 800 80368
rect 0 79432 800 79552
rect 139200 79296 140000 79416
rect 0 78616 800 78736
rect 0 77936 800 78056
rect 139200 78072 140000 78192
rect 0 77120 800 77240
rect 139200 76848 140000 76968
rect 0 76304 800 76424
rect 0 75624 800 75744
rect 139200 75488 140000 75608
rect 0 74808 800 74928
rect 139200 74264 140000 74384
rect 0 73992 800 74112
rect 0 73312 800 73432
rect 139200 73040 140000 73160
rect 0 72496 800 72616
rect 0 71680 800 71800
rect 139200 71680 140000 71800
rect 0 71000 800 71120
rect 139200 70456 140000 70576
rect 0 70184 800 70304
rect 0 69368 800 69488
rect 139200 69232 140000 69352
rect 0 68688 800 68808
rect 0 67872 800 67992
rect 139200 67872 140000 67992
rect 0 67056 800 67176
rect 139200 66648 140000 66768
rect 0 66376 800 66496
rect 0 65560 800 65680
rect 139200 65424 140000 65544
rect 0 64744 800 64864
rect 0 64064 800 64184
rect 139200 64064 140000 64184
rect 0 63248 800 63368
rect 139200 62840 140000 62960
rect 0 62432 800 62552
rect 0 61752 800 61872
rect 139200 61616 140000 61736
rect 0 60936 800 61056
rect 0 60256 800 60376
rect 139200 60256 140000 60376
rect 0 59440 800 59560
rect 139200 59032 140000 59152
rect 0 58624 800 58744
rect 0 57944 800 58064
rect 139200 57672 140000 57792
rect 0 57128 800 57248
rect 0 56312 800 56432
rect 139200 56448 140000 56568
rect 0 55632 800 55752
rect 139200 55224 140000 55344
rect 0 54816 800 54936
rect 0 54000 800 54120
rect 139200 53864 140000 53984
rect 0 53320 800 53440
rect 0 52504 800 52624
rect 139200 52640 140000 52760
rect 0 51688 800 51808
rect 139200 51416 140000 51536
rect 0 51008 800 51128
rect 0 50192 800 50312
rect 139200 50056 140000 50176
rect 0 49376 800 49496
rect 0 48696 800 48816
rect 139200 48832 140000 48952
rect 0 47880 800 48000
rect 139200 47608 140000 47728
rect 0 47064 800 47184
rect 0 46384 800 46504
rect 139200 46248 140000 46368
rect 0 45568 800 45688
rect 139200 45024 140000 45144
rect 0 44752 800 44872
rect 0 44072 800 44192
rect 139200 43800 140000 43920
rect 0 43256 800 43376
rect 0 42440 800 42560
rect 139200 42440 140000 42560
rect 0 41760 800 41880
rect 139200 41216 140000 41336
rect 0 40944 800 41064
rect 0 40264 800 40384
rect 139200 39856 140000 39976
rect 0 39448 800 39568
rect 0 38632 800 38752
rect 139200 38632 140000 38752
rect 0 37952 800 38072
rect 139200 37408 140000 37528
rect 0 37136 800 37256
rect 0 36320 800 36440
rect 139200 36048 140000 36168
rect 0 35640 800 35760
rect 0 34824 800 34944
rect 139200 34824 140000 34944
rect 0 34008 800 34128
rect 139200 33600 140000 33720
rect 0 33328 800 33448
rect 0 32512 800 32632
rect 139200 32240 140000 32360
rect 0 31696 800 31816
rect 0 31016 800 31136
rect 139200 31016 140000 31136
rect 0 30200 800 30320
rect 139200 29792 140000 29912
rect 0 29384 800 29504
rect 0 28704 800 28824
rect 139200 28432 140000 28552
rect 0 27888 800 28008
rect 0 27072 800 27192
rect 139200 27208 140000 27328
rect 0 26392 800 26512
rect 139200 25984 140000 26104
rect 0 25576 800 25696
rect 0 24760 800 24880
rect 139200 24624 140000 24744
rect 0 24080 800 24200
rect 0 23264 800 23384
rect 139200 23400 140000 23520
rect 0 22448 800 22568
rect 139200 22176 140000 22296
rect 0 21768 800 21888
rect 0 20952 800 21072
rect 139200 20816 140000 20936
rect 0 20272 800 20392
rect 0 19456 800 19576
rect 139200 19592 140000 19712
rect 0 18640 800 18760
rect 139200 18232 140000 18352
rect 0 17960 800 18080
rect 0 17144 800 17264
rect 139200 17008 140000 17128
rect 0 16328 800 16448
rect 0 15648 800 15768
rect 139200 15784 140000 15904
rect 0 14832 800 14952
rect 139200 14424 140000 14544
rect 0 14016 800 14136
rect 0 13336 800 13456
rect 139200 13200 140000 13320
rect 0 12520 800 12640
rect 139200 11976 140000 12096
rect 0 11704 800 11824
rect 0 11024 800 11144
rect 139200 10616 140000 10736
rect 0 10208 800 10328
rect 0 9392 800 9512
rect 139200 9392 140000 9512
rect 0 8712 800 8832
rect 139200 8168 140000 8288
rect 0 7896 800 8016
rect 0 7080 800 7200
rect 139200 6808 140000 6928
rect 0 6400 800 6520
rect 0 5584 800 5704
rect 139200 5584 140000 5704
rect 0 4768 800 4888
rect 139200 4360 140000 4480
rect 0 4088 800 4208
rect 0 3272 800 3392
rect 139200 3000 140000 3120
rect 0 2456 800 2576
rect 0 1776 800 1896
rect 139200 1776 140000 1896
rect 0 960 800 1080
rect 139200 552 140000 672
rect 0 280 800 400
<< obsm3 >>
rect 880 139336 139200 139501
rect 880 139328 139120 139336
rect 800 139056 139120 139328
rect 800 138792 139200 139056
rect 880 138512 139200 138792
rect 800 138112 139200 138512
rect 880 137832 139120 138112
rect 800 137296 139200 137832
rect 880 137016 139200 137296
rect 800 136752 139200 137016
rect 800 136480 139120 136752
rect 880 136472 139120 136480
rect 880 136200 139200 136472
rect 800 135800 139200 136200
rect 880 135528 139200 135800
rect 880 135520 139120 135528
rect 800 135248 139120 135520
rect 800 134984 139200 135248
rect 880 134704 139200 134984
rect 800 134304 139200 134704
rect 800 134168 139120 134304
rect 880 134024 139120 134168
rect 880 133888 139200 134024
rect 800 133488 139200 133888
rect 880 133208 139200 133488
rect 800 132944 139200 133208
rect 800 132672 139120 132944
rect 880 132664 139120 132672
rect 880 132392 139200 132664
rect 800 131856 139200 132392
rect 880 131720 139200 131856
rect 880 131576 139120 131720
rect 800 131440 139120 131576
rect 800 131176 139200 131440
rect 880 130896 139200 131176
rect 800 130496 139200 130896
rect 800 130360 139120 130496
rect 880 130216 139120 130360
rect 880 130080 139200 130216
rect 800 129544 139200 130080
rect 880 129264 139200 129544
rect 800 129136 139200 129264
rect 800 128864 139120 129136
rect 880 128856 139120 128864
rect 880 128584 139200 128856
rect 800 128048 139200 128584
rect 880 127912 139200 128048
rect 880 127768 139120 127912
rect 800 127632 139120 127768
rect 800 127232 139200 127632
rect 880 126952 139200 127232
rect 800 126688 139200 126952
rect 800 126552 139120 126688
rect 880 126408 139120 126552
rect 880 126272 139200 126408
rect 800 125736 139200 126272
rect 880 125456 139200 125736
rect 800 125328 139200 125456
rect 800 125048 139120 125328
rect 800 124920 139200 125048
rect 880 124640 139200 124920
rect 800 124240 139200 124640
rect 880 124104 139200 124240
rect 880 123960 139120 124104
rect 800 123824 139120 123960
rect 800 123424 139200 123824
rect 880 123144 139200 123424
rect 800 122880 139200 123144
rect 800 122608 139120 122880
rect 880 122600 139120 122608
rect 880 122328 139200 122600
rect 800 121928 139200 122328
rect 880 121648 139200 121928
rect 800 121520 139200 121648
rect 800 121240 139120 121520
rect 800 121112 139200 121240
rect 880 120832 139200 121112
rect 800 120432 139200 120832
rect 880 120296 139200 120432
rect 880 120152 139120 120296
rect 800 120016 139120 120152
rect 800 119616 139200 120016
rect 880 119336 139200 119616
rect 800 118936 139200 119336
rect 800 118800 139120 118936
rect 880 118656 139120 118800
rect 880 118520 139200 118656
rect 800 118120 139200 118520
rect 880 117840 139200 118120
rect 800 117712 139200 117840
rect 800 117432 139120 117712
rect 800 117304 139200 117432
rect 880 117024 139200 117304
rect 800 116488 139200 117024
rect 880 116208 139120 116488
rect 800 115808 139200 116208
rect 880 115528 139200 115808
rect 800 115128 139200 115528
rect 800 114992 139120 115128
rect 880 114848 139120 114992
rect 880 114712 139200 114848
rect 800 114176 139200 114712
rect 880 113904 139200 114176
rect 880 113896 139120 113904
rect 800 113624 139120 113896
rect 800 113496 139200 113624
rect 880 113216 139200 113496
rect 800 112680 139200 113216
rect 880 112400 139120 112680
rect 800 111864 139200 112400
rect 880 111584 139200 111864
rect 800 111320 139200 111584
rect 800 111184 139120 111320
rect 880 111040 139120 111184
rect 880 110904 139200 111040
rect 800 110368 139200 110904
rect 880 110096 139200 110368
rect 880 110088 139120 110096
rect 800 109816 139120 110088
rect 800 109552 139200 109816
rect 880 109272 139200 109552
rect 800 108872 139200 109272
rect 880 108592 139120 108872
rect 800 108056 139200 108592
rect 880 107776 139200 108056
rect 800 107512 139200 107776
rect 800 107240 139120 107512
rect 880 107232 139120 107240
rect 880 106960 139200 107232
rect 800 106560 139200 106960
rect 880 106288 139200 106560
rect 880 106280 139120 106288
rect 800 106008 139120 106280
rect 800 105744 139200 106008
rect 880 105464 139200 105744
rect 800 105064 139200 105464
rect 800 104928 139120 105064
rect 880 104784 139120 104928
rect 880 104648 139200 104784
rect 800 104248 139200 104648
rect 880 103968 139200 104248
rect 800 103704 139200 103968
rect 800 103432 139120 103704
rect 880 103424 139120 103432
rect 880 103152 139200 103424
rect 800 102616 139200 103152
rect 880 102480 139200 102616
rect 880 102336 139120 102480
rect 800 102200 139120 102336
rect 800 101936 139200 102200
rect 880 101656 139200 101936
rect 800 101256 139200 101656
rect 800 101120 139120 101256
rect 880 100976 139120 101120
rect 880 100840 139200 100976
rect 800 100440 139200 100840
rect 880 100160 139200 100440
rect 800 99896 139200 100160
rect 800 99624 139120 99896
rect 880 99616 139120 99624
rect 880 99344 139200 99616
rect 800 98808 139200 99344
rect 880 98672 139200 98808
rect 880 98528 139120 98672
rect 800 98392 139120 98528
rect 800 98128 139200 98392
rect 880 97848 139200 98128
rect 800 97312 139200 97848
rect 880 97032 139120 97312
rect 800 96496 139200 97032
rect 880 96216 139200 96496
rect 800 96088 139200 96216
rect 800 95816 139120 96088
rect 880 95808 139120 95816
rect 880 95536 139200 95808
rect 800 95000 139200 95536
rect 880 94864 139200 95000
rect 880 94720 139120 94864
rect 800 94584 139120 94720
rect 800 94184 139200 94584
rect 880 93904 139200 94184
rect 800 93504 139200 93904
rect 880 93224 139120 93504
rect 800 92688 139200 93224
rect 880 92408 139200 92688
rect 800 92280 139200 92408
rect 800 92000 139120 92280
rect 800 91872 139200 92000
rect 880 91592 139200 91872
rect 800 91192 139200 91592
rect 880 91056 139200 91192
rect 880 90912 139120 91056
rect 800 90776 139120 90912
rect 800 90376 139200 90776
rect 880 90096 139200 90376
rect 800 89696 139200 90096
rect 800 89560 139120 89696
rect 880 89416 139120 89560
rect 880 89280 139200 89416
rect 800 88880 139200 89280
rect 880 88600 139200 88880
rect 800 88472 139200 88600
rect 800 88192 139120 88472
rect 800 88064 139200 88192
rect 880 87784 139200 88064
rect 800 87248 139200 87784
rect 880 86968 139120 87248
rect 800 86568 139200 86968
rect 880 86288 139200 86568
rect 800 85888 139200 86288
rect 800 85752 139120 85888
rect 880 85608 139120 85752
rect 880 85472 139200 85608
rect 800 84936 139200 85472
rect 880 84664 139200 84936
rect 880 84656 139120 84664
rect 800 84384 139120 84656
rect 800 84256 139200 84384
rect 880 83976 139200 84256
rect 800 83440 139200 83976
rect 880 83160 139120 83440
rect 800 82624 139200 83160
rect 880 82344 139200 82624
rect 800 82080 139200 82344
rect 800 81944 139120 82080
rect 880 81800 139120 81944
rect 880 81664 139200 81800
rect 800 81128 139200 81664
rect 880 80856 139200 81128
rect 880 80848 139120 80856
rect 800 80576 139120 80848
rect 800 80448 139200 80576
rect 880 80168 139200 80448
rect 800 79632 139200 80168
rect 880 79496 139200 79632
rect 880 79352 139120 79496
rect 800 79216 139120 79352
rect 800 78816 139200 79216
rect 880 78536 139200 78816
rect 800 78272 139200 78536
rect 800 78136 139120 78272
rect 880 77992 139120 78136
rect 880 77856 139200 77992
rect 800 77320 139200 77856
rect 880 77048 139200 77320
rect 880 77040 139120 77048
rect 800 76768 139120 77040
rect 800 76504 139200 76768
rect 880 76224 139200 76504
rect 800 75824 139200 76224
rect 880 75688 139200 75824
rect 880 75544 139120 75688
rect 800 75408 139120 75544
rect 800 75008 139200 75408
rect 880 74728 139200 75008
rect 800 74464 139200 74728
rect 800 74192 139120 74464
rect 880 74184 139120 74192
rect 880 73912 139200 74184
rect 800 73512 139200 73912
rect 880 73240 139200 73512
rect 880 73232 139120 73240
rect 800 72960 139120 73232
rect 800 72696 139200 72960
rect 880 72416 139200 72696
rect 800 71880 139200 72416
rect 880 71600 139120 71880
rect 800 71200 139200 71600
rect 880 70920 139200 71200
rect 800 70656 139200 70920
rect 800 70384 139120 70656
rect 880 70376 139120 70384
rect 880 70104 139200 70376
rect 800 69568 139200 70104
rect 880 69432 139200 69568
rect 880 69288 139120 69432
rect 800 69152 139120 69288
rect 800 68888 139200 69152
rect 880 68608 139200 68888
rect 800 68072 139200 68608
rect 880 67792 139120 68072
rect 800 67256 139200 67792
rect 880 66976 139200 67256
rect 800 66848 139200 66976
rect 800 66576 139120 66848
rect 880 66568 139120 66576
rect 880 66296 139200 66568
rect 800 65760 139200 66296
rect 880 65624 139200 65760
rect 880 65480 139120 65624
rect 800 65344 139120 65480
rect 800 64944 139200 65344
rect 880 64664 139200 64944
rect 800 64264 139200 64664
rect 880 63984 139120 64264
rect 800 63448 139200 63984
rect 880 63168 139200 63448
rect 800 63040 139200 63168
rect 800 62760 139120 63040
rect 800 62632 139200 62760
rect 880 62352 139200 62632
rect 800 61952 139200 62352
rect 880 61816 139200 61952
rect 880 61672 139120 61816
rect 800 61536 139120 61672
rect 800 61136 139200 61536
rect 880 60856 139200 61136
rect 800 60456 139200 60856
rect 880 60176 139120 60456
rect 800 59640 139200 60176
rect 880 59360 139200 59640
rect 800 59232 139200 59360
rect 800 58952 139120 59232
rect 800 58824 139200 58952
rect 880 58544 139200 58824
rect 800 58144 139200 58544
rect 880 57872 139200 58144
rect 880 57864 139120 57872
rect 800 57592 139120 57864
rect 800 57328 139200 57592
rect 880 57048 139200 57328
rect 800 56648 139200 57048
rect 800 56512 139120 56648
rect 880 56368 139120 56512
rect 880 56232 139200 56368
rect 800 55832 139200 56232
rect 880 55552 139200 55832
rect 800 55424 139200 55552
rect 800 55144 139120 55424
rect 800 55016 139200 55144
rect 880 54736 139200 55016
rect 800 54200 139200 54736
rect 880 54064 139200 54200
rect 880 53920 139120 54064
rect 800 53784 139120 53920
rect 800 53520 139200 53784
rect 880 53240 139200 53520
rect 800 52840 139200 53240
rect 800 52704 139120 52840
rect 880 52560 139120 52704
rect 880 52424 139200 52560
rect 800 51888 139200 52424
rect 880 51616 139200 51888
rect 880 51608 139120 51616
rect 800 51336 139120 51608
rect 800 51208 139200 51336
rect 880 50928 139200 51208
rect 800 50392 139200 50928
rect 880 50256 139200 50392
rect 880 50112 139120 50256
rect 800 49976 139120 50112
rect 800 49576 139200 49976
rect 880 49296 139200 49576
rect 800 49032 139200 49296
rect 800 48896 139120 49032
rect 880 48752 139120 48896
rect 880 48616 139200 48752
rect 800 48080 139200 48616
rect 880 47808 139200 48080
rect 880 47800 139120 47808
rect 800 47528 139120 47800
rect 800 47264 139200 47528
rect 880 46984 139200 47264
rect 800 46584 139200 46984
rect 880 46448 139200 46584
rect 880 46304 139120 46448
rect 800 46168 139120 46304
rect 800 45768 139200 46168
rect 880 45488 139200 45768
rect 800 45224 139200 45488
rect 800 44952 139120 45224
rect 880 44944 139120 44952
rect 880 44672 139200 44944
rect 800 44272 139200 44672
rect 880 44000 139200 44272
rect 880 43992 139120 44000
rect 800 43720 139120 43992
rect 800 43456 139200 43720
rect 880 43176 139200 43456
rect 800 42640 139200 43176
rect 880 42360 139120 42640
rect 800 41960 139200 42360
rect 880 41680 139200 41960
rect 800 41416 139200 41680
rect 800 41144 139120 41416
rect 880 41136 139120 41144
rect 880 40864 139200 41136
rect 800 40464 139200 40864
rect 880 40184 139200 40464
rect 800 40056 139200 40184
rect 800 39776 139120 40056
rect 800 39648 139200 39776
rect 880 39368 139200 39648
rect 800 38832 139200 39368
rect 880 38552 139120 38832
rect 800 38152 139200 38552
rect 880 37872 139200 38152
rect 800 37608 139200 37872
rect 800 37336 139120 37608
rect 880 37328 139120 37336
rect 880 37056 139200 37328
rect 800 36520 139200 37056
rect 880 36248 139200 36520
rect 880 36240 139120 36248
rect 800 35968 139120 36240
rect 800 35840 139200 35968
rect 880 35560 139200 35840
rect 800 35024 139200 35560
rect 880 34744 139120 35024
rect 800 34208 139200 34744
rect 880 33928 139200 34208
rect 800 33800 139200 33928
rect 800 33528 139120 33800
rect 880 33520 139120 33528
rect 880 33248 139200 33520
rect 800 32712 139200 33248
rect 880 32440 139200 32712
rect 880 32432 139120 32440
rect 800 32160 139120 32432
rect 800 31896 139200 32160
rect 880 31616 139200 31896
rect 800 31216 139200 31616
rect 880 30936 139120 31216
rect 800 30400 139200 30936
rect 880 30120 139200 30400
rect 800 29992 139200 30120
rect 800 29712 139120 29992
rect 800 29584 139200 29712
rect 880 29304 139200 29584
rect 800 28904 139200 29304
rect 880 28632 139200 28904
rect 880 28624 139120 28632
rect 800 28352 139120 28624
rect 800 28088 139200 28352
rect 880 27808 139200 28088
rect 800 27408 139200 27808
rect 800 27272 139120 27408
rect 880 27128 139120 27272
rect 880 26992 139200 27128
rect 800 26592 139200 26992
rect 880 26312 139200 26592
rect 800 26184 139200 26312
rect 800 25904 139120 26184
rect 800 25776 139200 25904
rect 880 25496 139200 25776
rect 800 24960 139200 25496
rect 880 24824 139200 24960
rect 880 24680 139120 24824
rect 800 24544 139120 24680
rect 800 24280 139200 24544
rect 880 24000 139200 24280
rect 800 23600 139200 24000
rect 800 23464 139120 23600
rect 880 23320 139120 23464
rect 880 23184 139200 23320
rect 800 22648 139200 23184
rect 880 22376 139200 22648
rect 880 22368 139120 22376
rect 800 22096 139120 22368
rect 800 21968 139200 22096
rect 880 21688 139200 21968
rect 800 21152 139200 21688
rect 880 21016 139200 21152
rect 880 20872 139120 21016
rect 800 20736 139120 20872
rect 800 20472 139200 20736
rect 880 20192 139200 20472
rect 800 19792 139200 20192
rect 800 19656 139120 19792
rect 880 19512 139120 19656
rect 880 19376 139200 19512
rect 800 18840 139200 19376
rect 880 18560 139200 18840
rect 800 18432 139200 18560
rect 800 18160 139120 18432
rect 880 18152 139120 18160
rect 880 17880 139200 18152
rect 800 17344 139200 17880
rect 880 17208 139200 17344
rect 880 17064 139120 17208
rect 800 16928 139120 17064
rect 800 16528 139200 16928
rect 880 16248 139200 16528
rect 800 15984 139200 16248
rect 800 15848 139120 15984
rect 880 15704 139120 15848
rect 880 15568 139200 15704
rect 800 15032 139200 15568
rect 880 14752 139200 15032
rect 800 14624 139200 14752
rect 800 14344 139120 14624
rect 800 14216 139200 14344
rect 880 13936 139200 14216
rect 800 13536 139200 13936
rect 880 13400 139200 13536
rect 880 13256 139120 13400
rect 800 13120 139120 13256
rect 800 12720 139200 13120
rect 880 12440 139200 12720
rect 800 12176 139200 12440
rect 800 11904 139120 12176
rect 880 11896 139120 11904
rect 880 11624 139200 11896
rect 800 11224 139200 11624
rect 880 10944 139200 11224
rect 800 10816 139200 10944
rect 800 10536 139120 10816
rect 800 10408 139200 10536
rect 880 10128 139200 10408
rect 800 9592 139200 10128
rect 880 9312 139120 9592
rect 800 8912 139200 9312
rect 880 8632 139200 8912
rect 800 8368 139200 8632
rect 800 8096 139120 8368
rect 880 8088 139120 8096
rect 880 7816 139200 8088
rect 800 7280 139200 7816
rect 880 7008 139200 7280
rect 880 7000 139120 7008
rect 800 6728 139120 7000
rect 800 6600 139200 6728
rect 880 6320 139200 6600
rect 800 5784 139200 6320
rect 880 5504 139120 5784
rect 800 4968 139200 5504
rect 880 4688 139200 4968
rect 800 4560 139200 4688
rect 800 4288 139120 4560
rect 880 4280 139120 4288
rect 880 4008 139200 4280
rect 800 3472 139200 4008
rect 880 3200 139200 3472
rect 880 3192 139120 3200
rect 800 2920 139120 3192
rect 800 2656 139200 2920
rect 880 2376 139200 2656
rect 800 1976 139200 2376
rect 880 1696 139120 1976
rect 800 1160 139200 1696
rect 880 880 139200 1160
rect 800 752 139200 880
rect 800 480 139120 752
rect 880 472 139120 480
rect 880 307 139200 472
<< metal4 >>
rect 4208 2128 4528 137680
rect 19568 2128 19888 137680
rect 34928 2128 35248 137680
rect 50288 2128 50608 137680
rect 65648 2128 65968 137680
rect 81008 2128 81328 137680
rect 96368 2128 96688 137680
rect 111728 2128 112048 137680
rect 127088 2128 127408 137680
<< obsm4 >>
rect 2451 2347 4128 137189
rect 4608 2347 19488 137189
rect 19968 2347 34848 137189
rect 35328 2347 45021 137189
<< labels >>
rlabel metal2 s 3514 0 3570 800 6 clock
port 1 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 io_dbus_addr[0]
port 2 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 io_dbus_addr[10]
port 3 nsew signal input
rlabel metal3 s 0 31696 800 31816 6 io_dbus_addr[11]
port 4 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 io_dbus_addr[12]
port 5 nsew signal input
rlabel metal3 s 0 36320 800 36440 6 io_dbus_addr[13]
port 6 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 io_dbus_addr[14]
port 7 nsew signal input
rlabel metal3 s 0 40944 800 41064 6 io_dbus_addr[15]
port 8 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 io_dbus_addr[16]
port 9 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 io_dbus_addr[17]
port 10 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 io_dbus_addr[18]
port 11 nsew signal input
rlabel metal3 s 0 50192 800 50312 6 io_dbus_addr[19]
port 12 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 io_dbus_addr[1]
port 13 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 io_dbus_addr[20]
port 14 nsew signal input
rlabel metal3 s 0 54816 800 54936 6 io_dbus_addr[21]
port 15 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 io_dbus_addr[22]
port 16 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 io_dbus_addr[23]
port 17 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 io_dbus_addr[24]
port 18 nsew signal input
rlabel metal3 s 0 64064 800 64184 6 io_dbus_addr[25]
port 19 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 io_dbus_addr[26]
port 20 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 io_dbus_addr[27]
port 21 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 io_dbus_addr[28]
port 22 nsew signal input
rlabel metal3 s 0 73312 800 73432 6 io_dbus_addr[29]
port 23 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 io_dbus_addr[2]
port 24 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 io_dbus_addr[30]
port 25 nsew signal input
rlabel metal3 s 0 77936 800 78056 6 io_dbus_addr[31]
port 26 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 io_dbus_addr[3]
port 27 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 io_dbus_addr[4]
port 28 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 io_dbus_addr[5]
port 29 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 io_dbus_addr[6]
port 30 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 io_dbus_addr[7]
port 31 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 io_dbus_addr[8]
port 32 nsew signal input
rlabel metal3 s 0 27072 800 27192 6 io_dbus_addr[9]
port 33 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 io_dbus_ld_type[0]
port 34 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 io_dbus_ld_type[1]
port 35 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 io_dbus_ld_type[2]
port 36 nsew signal input
rlabel metal3 s 0 280 800 400 6 io_dbus_rd_en
port 37 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 io_dbus_rdata[0]
port 38 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 io_dbus_rdata[10]
port 39 nsew signal output
rlabel metal3 s 0 32512 800 32632 6 io_dbus_rdata[11]
port 40 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 io_dbus_rdata[12]
port 41 nsew signal output
rlabel metal3 s 0 37136 800 37256 6 io_dbus_rdata[13]
port 42 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 io_dbus_rdata[14]
port 43 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 io_dbus_rdata[15]
port 44 nsew signal output
rlabel metal3 s 0 44072 800 44192 6 io_dbus_rdata[16]
port 45 nsew signal output
rlabel metal3 s 0 46384 800 46504 6 io_dbus_rdata[17]
port 46 nsew signal output
rlabel metal3 s 0 48696 800 48816 6 io_dbus_rdata[18]
port 47 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 io_dbus_rdata[19]
port 48 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 io_dbus_rdata[1]
port 49 nsew signal output
rlabel metal3 s 0 53320 800 53440 6 io_dbus_rdata[20]
port 50 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 io_dbus_rdata[21]
port 51 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 io_dbus_rdata[22]
port 52 nsew signal output
rlabel metal3 s 0 60256 800 60376 6 io_dbus_rdata[23]
port 53 nsew signal output
rlabel metal3 s 0 62432 800 62552 6 io_dbus_rdata[24]
port 54 nsew signal output
rlabel metal3 s 0 64744 800 64864 6 io_dbus_rdata[25]
port 55 nsew signal output
rlabel metal3 s 0 67056 800 67176 6 io_dbus_rdata[26]
port 56 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 io_dbus_rdata[27]
port 57 nsew signal output
rlabel metal3 s 0 71680 800 71800 6 io_dbus_rdata[28]
port 58 nsew signal output
rlabel metal3 s 0 73992 800 74112 6 io_dbus_rdata[29]
port 59 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 io_dbus_rdata[2]
port 60 nsew signal output
rlabel metal3 s 0 76304 800 76424 6 io_dbus_rdata[30]
port 61 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 io_dbus_rdata[31]
port 62 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 io_dbus_rdata[3]
port 63 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 io_dbus_rdata[4]
port 64 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 io_dbus_rdata[5]
port 65 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 io_dbus_rdata[6]
port 66 nsew signal output
rlabel metal3 s 0 23264 800 23384 6 io_dbus_rdata[7]
port 67 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 io_dbus_rdata[8]
port 68 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 io_dbus_rdata[9]
port 69 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 io_dbus_st_type[0]
port 70 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 io_dbus_st_type[1]
port 71 nsew signal input
rlabel metal3 s 0 960 800 1080 6 io_dbus_valid
port 72 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 io_dbus_wdata[0]
port 73 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 io_dbus_wdata[10]
port 74 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 io_dbus_wdata[11]
port 75 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 io_dbus_wdata[12]
port 76 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 io_dbus_wdata[13]
port 77 nsew signal input
rlabel metal3 s 0 40264 800 40384 6 io_dbus_wdata[14]
port 78 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 io_dbus_wdata[15]
port 79 nsew signal input
rlabel metal3 s 0 44752 800 44872 6 io_dbus_wdata[16]
port 80 nsew signal input
rlabel metal3 s 0 47064 800 47184 6 io_dbus_wdata[17]
port 81 nsew signal input
rlabel metal3 s 0 49376 800 49496 6 io_dbus_wdata[18]
port 82 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 io_dbus_wdata[19]
port 83 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 io_dbus_wdata[1]
port 84 nsew signal input
rlabel metal3 s 0 54000 800 54120 6 io_dbus_wdata[20]
port 85 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 io_dbus_wdata[21]
port 86 nsew signal input
rlabel metal3 s 0 58624 800 58744 6 io_dbus_wdata[22]
port 87 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 io_dbus_wdata[23]
port 88 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 io_dbus_wdata[24]
port 89 nsew signal input
rlabel metal3 s 0 65560 800 65680 6 io_dbus_wdata[25]
port 90 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 io_dbus_wdata[26]
port 91 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 io_dbus_wdata[27]
port 92 nsew signal input
rlabel metal3 s 0 72496 800 72616 6 io_dbus_wdata[28]
port 93 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 io_dbus_wdata[29]
port 94 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 io_dbus_wdata[2]
port 95 nsew signal input
rlabel metal3 s 0 77120 800 77240 6 io_dbus_wdata[30]
port 96 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 io_dbus_wdata[31]
port 97 nsew signal input
rlabel metal3 s 0 14832 800 14952 6 io_dbus_wdata[3]
port 98 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 io_dbus_wdata[4]
port 99 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 io_dbus_wdata[5]
port 100 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 io_dbus_wdata[6]
port 101 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 io_dbus_wdata[7]
port 102 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 io_dbus_wdata[8]
port 103 nsew signal input
rlabel metal3 s 0 28704 800 28824 6 io_dbus_wdata[9]
port 104 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 io_dbus_wr_en
port 105 nsew signal input
rlabel metal2 s 3238 139200 3294 140000 6 io_dmem_io_addr[0]
port 106 nsew signal output
rlabel metal2 s 8390 139200 8446 140000 6 io_dmem_io_addr[1]
port 107 nsew signal output
rlabel metal2 s 13542 139200 13598 140000 6 io_dmem_io_addr[2]
port 108 nsew signal output
rlabel metal2 s 18786 139200 18842 140000 6 io_dmem_io_addr[3]
port 109 nsew signal output
rlabel metal2 s 23938 139200 23994 140000 6 io_dmem_io_addr[4]
port 110 nsew signal output
rlabel metal2 s 27802 139200 27858 140000 6 io_dmem_io_addr[5]
port 111 nsew signal output
rlabel metal2 s 31758 139200 31814 140000 6 io_dmem_io_addr[6]
port 112 nsew signal output
rlabel metal2 s 35622 139200 35678 140000 6 io_dmem_io_addr[7]
port 113 nsew signal output
rlabel metal2 s 662 139200 718 140000 6 io_dmem_io_cs
port 114 nsew signal output
rlabel metal2 s 4526 139200 4582 140000 6 io_dmem_io_rdata[0]
port 115 nsew signal input
rlabel metal2 s 44730 139200 44786 140000 6 io_dmem_io_rdata[10]
port 116 nsew signal input
rlabel metal2 s 47306 139200 47362 140000 6 io_dmem_io_rdata[11]
port 117 nsew signal input
rlabel metal2 s 49882 139200 49938 140000 6 io_dmem_io_rdata[12]
port 118 nsew signal input
rlabel metal2 s 52458 139200 52514 140000 6 io_dmem_io_rdata[13]
port 119 nsew signal input
rlabel metal2 s 55034 139200 55090 140000 6 io_dmem_io_rdata[14]
port 120 nsew signal input
rlabel metal2 s 57702 139200 57758 140000 6 io_dmem_io_rdata[15]
port 121 nsew signal input
rlabel metal2 s 60278 139200 60334 140000 6 io_dmem_io_rdata[16]
port 122 nsew signal input
rlabel metal2 s 62854 139200 62910 140000 6 io_dmem_io_rdata[17]
port 123 nsew signal input
rlabel metal2 s 65430 139200 65486 140000 6 io_dmem_io_rdata[18]
port 124 nsew signal input
rlabel metal2 s 68006 139200 68062 140000 6 io_dmem_io_rdata[19]
port 125 nsew signal input
rlabel metal2 s 9678 139200 9734 140000 6 io_dmem_io_rdata[1]
port 126 nsew signal input
rlabel metal2 s 70674 139200 70730 140000 6 io_dmem_io_rdata[20]
port 127 nsew signal input
rlabel metal2 s 73250 139200 73306 140000 6 io_dmem_io_rdata[21]
port 128 nsew signal input
rlabel metal2 s 75826 139200 75882 140000 6 io_dmem_io_rdata[22]
port 129 nsew signal input
rlabel metal2 s 78402 139200 78458 140000 6 io_dmem_io_rdata[23]
port 130 nsew signal input
rlabel metal2 s 80978 139200 81034 140000 6 io_dmem_io_rdata[24]
port 131 nsew signal input
rlabel metal2 s 83554 139200 83610 140000 6 io_dmem_io_rdata[25]
port 132 nsew signal input
rlabel metal2 s 86222 139200 86278 140000 6 io_dmem_io_rdata[26]
port 133 nsew signal input
rlabel metal2 s 88798 139200 88854 140000 6 io_dmem_io_rdata[27]
port 134 nsew signal input
rlabel metal2 s 91374 139200 91430 140000 6 io_dmem_io_rdata[28]
port 135 nsew signal input
rlabel metal2 s 93950 139200 94006 140000 6 io_dmem_io_rdata[29]
port 136 nsew signal input
rlabel metal2 s 14922 139200 14978 140000 6 io_dmem_io_rdata[2]
port 137 nsew signal input
rlabel metal2 s 96526 139200 96582 140000 6 io_dmem_io_rdata[30]
port 138 nsew signal input
rlabel metal2 s 99194 139200 99250 140000 6 io_dmem_io_rdata[31]
port 139 nsew signal input
rlabel metal2 s 20074 139200 20130 140000 6 io_dmem_io_rdata[3]
port 140 nsew signal input
rlabel metal2 s 25226 139200 25282 140000 6 io_dmem_io_rdata[4]
port 141 nsew signal input
rlabel metal2 s 29182 139200 29238 140000 6 io_dmem_io_rdata[5]
port 142 nsew signal input
rlabel metal2 s 33046 139200 33102 140000 6 io_dmem_io_rdata[6]
port 143 nsew signal input
rlabel metal2 s 36910 139200 36966 140000 6 io_dmem_io_rdata[7]
port 144 nsew signal input
rlabel metal2 s 39486 139200 39542 140000 6 io_dmem_io_rdata[8]
port 145 nsew signal input
rlabel metal2 s 42062 139200 42118 140000 6 io_dmem_io_rdata[9]
port 146 nsew signal input
rlabel metal2 s 5814 139200 5870 140000 6 io_dmem_io_st_type[0]
port 147 nsew signal output
rlabel metal2 s 10966 139200 11022 140000 6 io_dmem_io_st_type[1]
port 148 nsew signal output
rlabel metal2 s 16210 139200 16266 140000 6 io_dmem_io_st_type[2]
port 149 nsew signal output
rlabel metal2 s 21362 139200 21418 140000 6 io_dmem_io_st_type[3]
port 150 nsew signal output
rlabel metal2 s 7102 139200 7158 140000 6 io_dmem_io_wdata[0]
port 151 nsew signal output
rlabel metal2 s 46018 139200 46074 140000 6 io_dmem_io_wdata[10]
port 152 nsew signal output
rlabel metal2 s 48594 139200 48650 140000 6 io_dmem_io_wdata[11]
port 153 nsew signal output
rlabel metal2 s 51170 139200 51226 140000 6 io_dmem_io_wdata[12]
port 154 nsew signal output
rlabel metal2 s 53746 139200 53802 140000 6 io_dmem_io_wdata[13]
port 155 nsew signal output
rlabel metal2 s 56322 139200 56378 140000 6 io_dmem_io_wdata[14]
port 156 nsew signal output
rlabel metal2 s 58990 139200 59046 140000 6 io_dmem_io_wdata[15]
port 157 nsew signal output
rlabel metal2 s 61566 139200 61622 140000 6 io_dmem_io_wdata[16]
port 158 nsew signal output
rlabel metal2 s 64142 139200 64198 140000 6 io_dmem_io_wdata[17]
port 159 nsew signal output
rlabel metal2 s 66718 139200 66774 140000 6 io_dmem_io_wdata[18]
port 160 nsew signal output
rlabel metal2 s 69294 139200 69350 140000 6 io_dmem_io_wdata[19]
port 161 nsew signal output
rlabel metal2 s 12254 139200 12310 140000 6 io_dmem_io_wdata[1]
port 162 nsew signal output
rlabel metal2 s 71962 139200 72018 140000 6 io_dmem_io_wdata[20]
port 163 nsew signal output
rlabel metal2 s 74538 139200 74594 140000 6 io_dmem_io_wdata[21]
port 164 nsew signal output
rlabel metal2 s 77114 139200 77170 140000 6 io_dmem_io_wdata[22]
port 165 nsew signal output
rlabel metal2 s 79690 139200 79746 140000 6 io_dmem_io_wdata[23]
port 166 nsew signal output
rlabel metal2 s 82266 139200 82322 140000 6 io_dmem_io_wdata[24]
port 167 nsew signal output
rlabel metal2 s 84934 139200 84990 140000 6 io_dmem_io_wdata[25]
port 168 nsew signal output
rlabel metal2 s 87510 139200 87566 140000 6 io_dmem_io_wdata[26]
port 169 nsew signal output
rlabel metal2 s 90086 139200 90142 140000 6 io_dmem_io_wdata[27]
port 170 nsew signal output
rlabel metal2 s 92662 139200 92718 140000 6 io_dmem_io_wdata[28]
port 171 nsew signal output
rlabel metal2 s 95238 139200 95294 140000 6 io_dmem_io_wdata[29]
port 172 nsew signal output
rlabel metal2 s 17498 139200 17554 140000 6 io_dmem_io_wdata[2]
port 173 nsew signal output
rlabel metal2 s 97814 139200 97870 140000 6 io_dmem_io_wdata[30]
port 174 nsew signal output
rlabel metal2 s 100482 139200 100538 140000 6 io_dmem_io_wdata[31]
port 175 nsew signal output
rlabel metal2 s 22650 139200 22706 140000 6 io_dmem_io_wdata[3]
port 176 nsew signal output
rlabel metal2 s 26514 139200 26570 140000 6 io_dmem_io_wdata[4]
port 177 nsew signal output
rlabel metal2 s 30470 139200 30526 140000 6 io_dmem_io_wdata[5]
port 178 nsew signal output
rlabel metal2 s 34334 139200 34390 140000 6 io_dmem_io_wdata[6]
port 179 nsew signal output
rlabel metal2 s 38198 139200 38254 140000 6 io_dmem_io_wdata[7]
port 180 nsew signal output
rlabel metal2 s 40774 139200 40830 140000 6 io_dmem_io_wdata[8]
port 181 nsew signal output
rlabel metal2 s 43442 139200 43498 140000 6 io_dmem_io_wdata[9]
port 182 nsew signal output
rlabel metal2 s 1950 139200 2006 140000 6 io_dmem_io_wr_en
port 183 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 io_ibus_addr[0]
port 184 nsew signal input
rlabel metal3 s 0 96296 800 96416 6 io_ibus_addr[10]
port 185 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 io_ibus_addr[11]
port 186 nsew signal input
rlabel metal3 s 0 99424 800 99544 6 io_ibus_addr[12]
port 187 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 io_ibus_addr[13]
port 188 nsew signal input
rlabel metal3 s 0 102416 800 102536 6 io_ibus_addr[14]
port 189 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 io_ibus_addr[15]
port 190 nsew signal input
rlabel metal3 s 0 105544 800 105664 6 io_ibus_addr[16]
port 191 nsew signal input
rlabel metal3 s 0 107040 800 107160 6 io_ibus_addr[17]
port 192 nsew signal input
rlabel metal3 s 0 108672 800 108792 6 io_ibus_addr[18]
port 193 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 io_ibus_addr[19]
port 194 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 io_ibus_addr[1]
port 195 nsew signal input
rlabel metal3 s 0 111664 800 111784 6 io_ibus_addr[20]
port 196 nsew signal input
rlabel metal3 s 0 113296 800 113416 6 io_ibus_addr[21]
port 197 nsew signal input
rlabel metal3 s 0 114792 800 114912 6 io_ibus_addr[22]
port 198 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 io_ibus_addr[23]
port 199 nsew signal input
rlabel metal3 s 0 117920 800 118040 6 io_ibus_addr[24]
port 200 nsew signal input
rlabel metal3 s 0 119416 800 119536 6 io_ibus_addr[25]
port 201 nsew signal input
rlabel metal3 s 0 120912 800 121032 6 io_ibus_addr[26]
port 202 nsew signal input
rlabel metal3 s 0 122408 800 122528 6 io_ibus_addr[27]
port 203 nsew signal input
rlabel metal3 s 0 124040 800 124160 6 io_ibus_addr[28]
port 204 nsew signal input
rlabel metal3 s 0 125536 800 125656 6 io_ibus_addr[29]
port 205 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 io_ibus_addr[2]
port 206 nsew signal input
rlabel metal3 s 0 127032 800 127152 6 io_ibus_addr[30]
port 207 nsew signal input
rlabel metal3 s 0 128664 800 128784 6 io_ibus_addr[31]
port 208 nsew signal input
rlabel metal3 s 0 85552 800 85672 6 io_ibus_addr[3]
port 209 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 io_ibus_addr[4]
port 210 nsew signal input
rlabel metal3 s 0 88680 800 88800 6 io_ibus_addr[5]
port 211 nsew signal input
rlabel metal3 s 0 90176 800 90296 6 io_ibus_addr[6]
port 212 nsew signal input
rlabel metal3 s 0 91672 800 91792 6 io_ibus_addr[7]
port 213 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 io_ibus_addr[8]
port 214 nsew signal input
rlabel metal3 s 0 94800 800 94920 6 io_ibus_addr[9]
port 215 nsew signal input
rlabel metal3 s 0 81744 800 81864 6 io_ibus_inst[0]
port 216 nsew signal output
rlabel metal3 s 0 97112 800 97232 6 io_ibus_inst[10]
port 217 nsew signal output
rlabel metal3 s 0 98608 800 98728 6 io_ibus_inst[11]
port 218 nsew signal output
rlabel metal3 s 0 100240 800 100360 6 io_ibus_inst[12]
port 219 nsew signal output
rlabel metal3 s 0 101736 800 101856 6 io_ibus_inst[13]
port 220 nsew signal output
rlabel metal3 s 0 103232 800 103352 6 io_ibus_inst[14]
port 221 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 io_ibus_inst[15]
port 222 nsew signal output
rlabel metal3 s 0 106360 800 106480 6 io_ibus_inst[16]
port 223 nsew signal output
rlabel metal3 s 0 107856 800 107976 6 io_ibus_inst[17]
port 224 nsew signal output
rlabel metal3 s 0 109352 800 109472 6 io_ibus_inst[18]
port 225 nsew signal output
rlabel metal3 s 0 110984 800 111104 6 io_ibus_inst[19]
port 226 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 io_ibus_inst[1]
port 227 nsew signal output
rlabel metal3 s 0 112480 800 112600 6 io_ibus_inst[20]
port 228 nsew signal output
rlabel metal3 s 0 113976 800 114096 6 io_ibus_inst[21]
port 229 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 io_ibus_inst[22]
port 230 nsew signal output
rlabel metal3 s 0 117104 800 117224 6 io_ibus_inst[23]
port 231 nsew signal output
rlabel metal3 s 0 118600 800 118720 6 io_ibus_inst[24]
port 232 nsew signal output
rlabel metal3 s 0 120232 800 120352 6 io_ibus_inst[25]
port 233 nsew signal output
rlabel metal3 s 0 121728 800 121848 6 io_ibus_inst[26]
port 234 nsew signal output
rlabel metal3 s 0 123224 800 123344 6 io_ibus_inst[27]
port 235 nsew signal output
rlabel metal3 s 0 124720 800 124840 6 io_ibus_inst[28]
port 236 nsew signal output
rlabel metal3 s 0 126352 800 126472 6 io_ibus_inst[29]
port 237 nsew signal output
rlabel metal3 s 0 84736 800 84856 6 io_ibus_inst[2]
port 238 nsew signal output
rlabel metal3 s 0 127848 800 127968 6 io_ibus_inst[30]
port 239 nsew signal output
rlabel metal3 s 0 129344 800 129464 6 io_ibus_inst[31]
port 240 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 io_ibus_inst[3]
port 241 nsew signal output
rlabel metal3 s 0 87864 800 87984 6 io_ibus_inst[4]
port 242 nsew signal output
rlabel metal3 s 0 89360 800 89480 6 io_ibus_inst[5]
port 243 nsew signal output
rlabel metal3 s 0 90992 800 91112 6 io_ibus_inst[6]
port 244 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 io_ibus_inst[7]
port 245 nsew signal output
rlabel metal3 s 0 93984 800 94104 6 io_ibus_inst[8]
port 246 nsew signal output
rlabel metal3 s 0 95616 800 95736 6 io_ibus_inst[9]
port 247 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 io_ibus_valid
port 248 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 io_imem_io_addr[0]
port 249 nsew signal output
rlabel metal2 s 103058 139200 103114 140000 6 io_imem_io_addr[1]
port 250 nsew signal output
rlabel metal2 s 104346 139200 104402 140000 6 io_imem_io_addr[2]
port 251 nsew signal output
rlabel metal3 s 139200 121320 140000 121440 6 io_imem_io_addr[3]
port 252 nsew signal output
rlabel metal2 s 108210 139200 108266 140000 6 io_imem_io_addr[4]
port 253 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 io_imem_io_addr[5]
port 254 nsew signal output
rlabel metal2 s 112074 139200 112130 140000 6 io_imem_io_addr[6]
port 255 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 io_imem_io_addr[7]
port 256 nsew signal output
rlabel metal3 s 0 133968 800 134088 6 io_imem_io_addr[8]
port 257 nsew signal output
rlabel metal3 s 139200 117512 140000 117632 6 io_imem_io_cs
port 258 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 io_imem_io_rdata[0]
port 259 nsew signal input
rlabel metal3 s 139200 128936 140000 129056 6 io_imem_io_rdata[10]
port 260 nsew signal input
rlabel metal2 s 114742 139200 114798 140000 6 io_imem_io_rdata[11]
port 261 nsew signal input
rlabel metal2 s 116030 139200 116086 140000 6 io_imem_io_rdata[12]
port 262 nsew signal input
rlabel metal2 s 117318 139200 117374 140000 6 io_imem_io_rdata[13]
port 263 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 io_imem_io_rdata[14]
port 264 nsew signal input
rlabel metal2 s 119894 139200 119950 140000 6 io_imem_io_rdata[15]
port 265 nsew signal input
rlabel metal2 s 122470 139200 122526 140000 6 io_imem_io_rdata[16]
port 266 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 io_imem_io_rdata[17]
port 267 nsew signal input
rlabel metal3 s 139200 134104 140000 134224 6 io_imem_io_rdata[18]
port 268 nsew signal input
rlabel metal2 s 123758 139200 123814 140000 6 io_imem_io_rdata[19]
port 269 nsew signal input
rlabel metal3 s 139200 118736 140000 118856 6 io_imem_io_rdata[1]
port 270 nsew signal input
rlabel metal3 s 139200 136552 140000 136672 6 io_imem_io_rdata[20]
port 271 nsew signal input
rlabel metal2 s 126334 139200 126390 140000 6 io_imem_io_rdata[21]
port 272 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 io_imem_io_rdata[22]
port 273 nsew signal input
rlabel metal3 s 139200 137912 140000 138032 6 io_imem_io_rdata[23]
port 274 nsew signal input
rlabel metal2 s 131578 139200 131634 140000 6 io_imem_io_rdata[24]
port 275 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 io_imem_io_rdata[25]
port 276 nsew signal input
rlabel metal3 s 0 138592 800 138712 6 io_imem_io_rdata[26]
port 277 nsew signal input
rlabel metal3 s 139200 139136 140000 139256 6 io_imem_io_rdata[27]
port 278 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 io_imem_io_rdata[28]
port 279 nsew signal input
rlabel metal2 s 135442 139200 135498 140000 6 io_imem_io_rdata[29]
port 280 nsew signal input
rlabel metal2 s 105634 139200 105690 140000 6 io_imem_io_rdata[2]
port 281 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 io_imem_io_rdata[30]
port 282 nsew signal input
rlabel metal2 s 139306 139200 139362 140000 6 io_imem_io_rdata[31]
port 283 nsew signal input
rlabel metal3 s 0 132472 800 132592 6 io_imem_io_rdata[3]
port 284 nsew signal input
rlabel metal2 s 109498 139200 109554 140000 6 io_imem_io_rdata[4]
port 285 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 io_imem_io_rdata[5]
port 286 nsew signal input
rlabel metal3 s 139200 125128 140000 125248 6 io_imem_io_rdata[6]
port 287 nsew signal input
rlabel metal3 s 139200 126488 140000 126608 6 io_imem_io_rdata[7]
port 288 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 io_imem_io_rdata[8]
port 289 nsew signal input
rlabel metal2 s 113454 139200 113510 140000 6 io_imem_io_rdata[9]
port 290 nsew signal input
rlabel metal3 s 0 131656 800 131776 6 io_imem_io_wdata[0]
port 291 nsew signal output
rlabel metal3 s 139200 130296 140000 130416 6 io_imem_io_wdata[10]
port 292 nsew signal output
rlabel metal3 s 0 135600 800 135720 6 io_imem_io_wdata[11]
port 293 nsew signal output
rlabel metal3 s 139200 131520 140000 131640 6 io_imem_io_wdata[12]
port 294 nsew signal output
rlabel metal2 s 118606 139200 118662 140000 6 io_imem_io_wdata[13]
port 295 nsew signal output
rlabel metal3 s 139200 132744 140000 132864 6 io_imem_io_wdata[14]
port 296 nsew signal output
rlabel metal2 s 121182 139200 121238 140000 6 io_imem_io_wdata[15]
port 297 nsew signal output
rlabel metal3 s 0 136280 800 136400 6 io_imem_io_wdata[16]
port 298 nsew signal output
rlabel metal3 s 0 137096 800 137216 6 io_imem_io_wdata[17]
port 299 nsew signal output
rlabel metal3 s 139200 135328 140000 135448 6 io_imem_io_wdata[18]
port 300 nsew signal output
rlabel metal3 s 0 137912 800 138032 6 io_imem_io_wdata[19]
port 301 nsew signal output
rlabel metal3 s 139200 120096 140000 120216 6 io_imem_io_wdata[1]
port 302 nsew signal output
rlabel metal2 s 125046 139200 125102 140000 6 io_imem_io_wdata[20]
port 303 nsew signal output
rlabel metal2 s 127714 139200 127770 140000 6 io_imem_io_wdata[21]
port 304 nsew signal output
rlabel metal2 s 129002 139200 129058 140000 6 io_imem_io_wdata[22]
port 305 nsew signal output
rlabel metal2 s 130290 139200 130346 140000 6 io_imem_io_wdata[23]
port 306 nsew signal output
rlabel metal2 s 132866 139200 132922 140000 6 io_imem_io_wdata[24]
port 307 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 io_imem_io_wdata[25]
port 308 nsew signal output
rlabel metal2 s 134154 139200 134210 140000 6 io_imem_io_wdata[26]
port 309 nsew signal output
rlabel metal3 s 0 139408 800 139528 6 io_imem_io_wdata[27]
port 310 nsew signal output
rlabel metal2 s 122470 0 122526 800 6 io_imem_io_wdata[28]
port 311 nsew signal output
rlabel metal2 s 136730 139200 136786 140000 6 io_imem_io_wdata[29]
port 312 nsew signal output
rlabel metal2 s 106922 139200 106978 140000 6 io_imem_io_wdata[2]
port 313 nsew signal output
rlabel metal2 s 138018 139200 138074 140000 6 io_imem_io_wdata[30]
port 314 nsew signal output
rlabel metal2 s 136454 0 136510 800 6 io_imem_io_wdata[31]
port 315 nsew signal output
rlabel metal3 s 139200 122680 140000 122800 6 io_imem_io_wdata[3]
port 316 nsew signal output
rlabel metal3 s 139200 123904 140000 124024 6 io_imem_io_wdata[4]
port 317 nsew signal output
rlabel metal2 s 110786 139200 110842 140000 6 io_imem_io_wdata[5]
port 318 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 io_imem_io_wdata[6]
port 319 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 io_imem_io_wdata[7]
port 320 nsew signal output
rlabel metal3 s 139200 127712 140000 127832 6 io_imem_io_wdata[8]
port 321 nsew signal output
rlabel metal3 s 0 134784 800 134904 6 io_imem_io_wdata[9]
port 322 nsew signal output
rlabel metal2 s 101770 139200 101826 140000 6 io_imem_io_wr_en
port 323 nsew signal output
rlabel metal3 s 139200 552 140000 672 6 io_motor_ack_i
port 324 nsew signal input
rlabel metal3 s 139200 1776 140000 1896 6 io_motor_addr_sel
port 325 nsew signal output
rlabel metal3 s 139200 3000 140000 3120 6 io_motor_data_i[0]
port 326 nsew signal input
rlabel metal3 s 139200 15784 140000 15904 6 io_motor_data_i[10]
port 327 nsew signal input
rlabel metal3 s 139200 17008 140000 17128 6 io_motor_data_i[11]
port 328 nsew signal input
rlabel metal3 s 139200 18232 140000 18352 6 io_motor_data_i[12]
port 329 nsew signal input
rlabel metal3 s 139200 19592 140000 19712 6 io_motor_data_i[13]
port 330 nsew signal input
rlabel metal3 s 139200 20816 140000 20936 6 io_motor_data_i[14]
port 331 nsew signal input
rlabel metal3 s 139200 22176 140000 22296 6 io_motor_data_i[15]
port 332 nsew signal input
rlabel metal3 s 139200 23400 140000 23520 6 io_motor_data_i[16]
port 333 nsew signal input
rlabel metal3 s 139200 24624 140000 24744 6 io_motor_data_i[17]
port 334 nsew signal input
rlabel metal3 s 139200 25984 140000 26104 6 io_motor_data_i[18]
port 335 nsew signal input
rlabel metal3 s 139200 27208 140000 27328 6 io_motor_data_i[19]
port 336 nsew signal input
rlabel metal3 s 139200 4360 140000 4480 6 io_motor_data_i[1]
port 337 nsew signal input
rlabel metal3 s 139200 28432 140000 28552 6 io_motor_data_i[20]
port 338 nsew signal input
rlabel metal3 s 139200 29792 140000 29912 6 io_motor_data_i[21]
port 339 nsew signal input
rlabel metal3 s 139200 31016 140000 31136 6 io_motor_data_i[22]
port 340 nsew signal input
rlabel metal3 s 139200 32240 140000 32360 6 io_motor_data_i[23]
port 341 nsew signal input
rlabel metal3 s 139200 33600 140000 33720 6 io_motor_data_i[24]
port 342 nsew signal input
rlabel metal3 s 139200 34824 140000 34944 6 io_motor_data_i[25]
port 343 nsew signal input
rlabel metal3 s 139200 36048 140000 36168 6 io_motor_data_i[26]
port 344 nsew signal input
rlabel metal3 s 139200 37408 140000 37528 6 io_motor_data_i[27]
port 345 nsew signal input
rlabel metal3 s 139200 38632 140000 38752 6 io_motor_data_i[28]
port 346 nsew signal input
rlabel metal3 s 139200 39856 140000 39976 6 io_motor_data_i[29]
port 347 nsew signal input
rlabel metal3 s 139200 5584 140000 5704 6 io_motor_data_i[2]
port 348 nsew signal input
rlabel metal3 s 139200 41216 140000 41336 6 io_motor_data_i[30]
port 349 nsew signal input
rlabel metal3 s 139200 42440 140000 42560 6 io_motor_data_i[31]
port 350 nsew signal input
rlabel metal3 s 139200 6808 140000 6928 6 io_motor_data_i[3]
port 351 nsew signal input
rlabel metal3 s 139200 8168 140000 8288 6 io_motor_data_i[4]
port 352 nsew signal input
rlabel metal3 s 139200 9392 140000 9512 6 io_motor_data_i[5]
port 353 nsew signal input
rlabel metal3 s 139200 10616 140000 10736 6 io_motor_data_i[6]
port 354 nsew signal input
rlabel metal3 s 139200 11976 140000 12096 6 io_motor_data_i[7]
port 355 nsew signal input
rlabel metal3 s 139200 13200 140000 13320 6 io_motor_data_i[8]
port 356 nsew signal input
rlabel metal3 s 139200 14424 140000 14544 6 io_motor_data_i[9]
port 357 nsew signal input
rlabel metal3 s 139200 112480 140000 112600 6 io_spi_clk
port 358 nsew signal output
rlabel metal3 s 139200 113704 140000 113824 6 io_spi_cs
port 359 nsew signal output
rlabel metal3 s 0 130160 800 130280 6 io_spi_irq
port 360 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 io_spi_miso
port 361 nsew signal input
rlabel metal3 s 139200 114928 140000 115048 6 io_spi_mosi
port 362 nsew signal output
rlabel metal3 s 0 130976 800 131096 6 io_uart_irq
port 363 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 io_uart_rx
port 364 nsew signal input
rlabel metal3 s 139200 116288 140000 116408 6 io_uart_tx
port 365 nsew signal output
rlabel metal3 s 139200 46248 140000 46368 6 io_wbm_m2s_addr[0]
port 366 nsew signal output
rlabel metal3 s 139200 76848 140000 76968 6 io_wbm_m2s_addr[10]
port 367 nsew signal output
rlabel metal3 s 139200 79296 140000 79416 6 io_wbm_m2s_addr[11]
port 368 nsew signal output
rlabel metal3 s 139200 81880 140000 82000 6 io_wbm_m2s_addr[12]
port 369 nsew signal output
rlabel metal3 s 139200 84464 140000 84584 6 io_wbm_m2s_addr[13]
port 370 nsew signal output
rlabel metal3 s 139200 87048 140000 87168 6 io_wbm_m2s_addr[14]
port 371 nsew signal output
rlabel metal3 s 139200 89496 140000 89616 6 io_wbm_m2s_addr[15]
port 372 nsew signal output
rlabel metal3 s 139200 50056 140000 50176 6 io_wbm_m2s_addr[1]
port 373 nsew signal output
rlabel metal3 s 139200 53864 140000 53984 6 io_wbm_m2s_addr[2]
port 374 nsew signal output
rlabel metal3 s 139200 57672 140000 57792 6 io_wbm_m2s_addr[3]
port 375 nsew signal output
rlabel metal3 s 139200 61616 140000 61736 6 io_wbm_m2s_addr[4]
port 376 nsew signal output
rlabel metal3 s 139200 64064 140000 64184 6 io_wbm_m2s_addr[5]
port 377 nsew signal output
rlabel metal3 s 139200 66648 140000 66768 6 io_wbm_m2s_addr[6]
port 378 nsew signal output
rlabel metal3 s 139200 69232 140000 69352 6 io_wbm_m2s_addr[7]
port 379 nsew signal output
rlabel metal3 s 139200 71680 140000 71800 6 io_wbm_m2s_addr[8]
port 380 nsew signal output
rlabel metal3 s 139200 74264 140000 74384 6 io_wbm_m2s_addr[9]
port 381 nsew signal output
rlabel metal3 s 139200 47608 140000 47728 6 io_wbm_m2s_data[0]
port 382 nsew signal output
rlabel metal3 s 139200 78072 140000 78192 6 io_wbm_m2s_data[10]
port 383 nsew signal output
rlabel metal3 s 139200 80656 140000 80776 6 io_wbm_m2s_data[11]
port 384 nsew signal output
rlabel metal3 s 139200 83240 140000 83360 6 io_wbm_m2s_data[12]
port 385 nsew signal output
rlabel metal3 s 139200 85688 140000 85808 6 io_wbm_m2s_data[13]
port 386 nsew signal output
rlabel metal3 s 139200 88272 140000 88392 6 io_wbm_m2s_data[14]
port 387 nsew signal output
rlabel metal3 s 139200 90856 140000 90976 6 io_wbm_m2s_data[15]
port 388 nsew signal output
rlabel metal3 s 139200 92080 140000 92200 6 io_wbm_m2s_data[16]
port 389 nsew signal output
rlabel metal3 s 139200 93304 140000 93424 6 io_wbm_m2s_data[17]
port 390 nsew signal output
rlabel metal3 s 139200 94664 140000 94784 6 io_wbm_m2s_data[18]
port 391 nsew signal output
rlabel metal3 s 139200 95888 140000 96008 6 io_wbm_m2s_data[19]
port 392 nsew signal output
rlabel metal3 s 139200 51416 140000 51536 6 io_wbm_m2s_data[1]
port 393 nsew signal output
rlabel metal3 s 139200 97112 140000 97232 6 io_wbm_m2s_data[20]
port 394 nsew signal output
rlabel metal3 s 139200 98472 140000 98592 6 io_wbm_m2s_data[21]
port 395 nsew signal output
rlabel metal3 s 139200 99696 140000 99816 6 io_wbm_m2s_data[22]
port 396 nsew signal output
rlabel metal3 s 139200 101056 140000 101176 6 io_wbm_m2s_data[23]
port 397 nsew signal output
rlabel metal3 s 139200 102280 140000 102400 6 io_wbm_m2s_data[24]
port 398 nsew signal output
rlabel metal3 s 139200 103504 140000 103624 6 io_wbm_m2s_data[25]
port 399 nsew signal output
rlabel metal3 s 139200 104864 140000 104984 6 io_wbm_m2s_data[26]
port 400 nsew signal output
rlabel metal3 s 139200 106088 140000 106208 6 io_wbm_m2s_data[27]
port 401 nsew signal output
rlabel metal3 s 139200 107312 140000 107432 6 io_wbm_m2s_data[28]
port 402 nsew signal output
rlabel metal3 s 139200 108672 140000 108792 6 io_wbm_m2s_data[29]
port 403 nsew signal output
rlabel metal3 s 139200 55224 140000 55344 6 io_wbm_m2s_data[2]
port 404 nsew signal output
rlabel metal3 s 139200 109896 140000 110016 6 io_wbm_m2s_data[30]
port 405 nsew signal output
rlabel metal3 s 139200 111120 140000 111240 6 io_wbm_m2s_data[31]
port 406 nsew signal output
rlabel metal3 s 139200 59032 140000 59152 6 io_wbm_m2s_data[3]
port 407 nsew signal output
rlabel metal3 s 139200 62840 140000 62960 6 io_wbm_m2s_data[4]
port 408 nsew signal output
rlabel metal3 s 139200 65424 140000 65544 6 io_wbm_m2s_data[5]
port 409 nsew signal output
rlabel metal3 s 139200 67872 140000 67992 6 io_wbm_m2s_data[6]
port 410 nsew signal output
rlabel metal3 s 139200 70456 140000 70576 6 io_wbm_m2s_data[7]
port 411 nsew signal output
rlabel metal3 s 139200 73040 140000 73160 6 io_wbm_m2s_data[8]
port 412 nsew signal output
rlabel metal3 s 139200 75488 140000 75608 6 io_wbm_m2s_data[9]
port 413 nsew signal output
rlabel metal3 s 139200 48832 140000 48952 6 io_wbm_m2s_sel[0]
port 414 nsew signal output
rlabel metal3 s 139200 52640 140000 52760 6 io_wbm_m2s_sel[1]
port 415 nsew signal output
rlabel metal3 s 139200 56448 140000 56568 6 io_wbm_m2s_sel[2]
port 416 nsew signal output
rlabel metal3 s 139200 60256 140000 60376 6 io_wbm_m2s_sel[3]
port 417 nsew signal output
rlabel metal3 s 139200 43800 140000 43920 6 io_wbm_m2s_stb
port 418 nsew signal output
rlabel metal3 s 139200 45024 140000 45144 6 io_wbm_m2s_we
port 419 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 reset
port 420 nsew signal input
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 421 nsew power input
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 421 nsew power input
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 421 nsew power input
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 421 nsew power input
rlabel metal4 s 127088 2128 127408 137680 6 vccd1
port 421 nsew power input
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 422 nsew ground input
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 422 nsew ground input
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 422 nsew ground input
rlabel metal4 s 111728 2128 112048 137680 6 vssd1
port 422 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 140000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11497784
string GDS_FILE /home/em/mpw/UETRV-ECORE/openlane/Wishbone_InterConnect/runs/Wishbone_InterConnect/results/finishing/WB_InterConnect.magic.gds
string GDS_START 903408
<< end >>

