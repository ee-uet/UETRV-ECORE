module IMem_Interface( // @[:@3093.2]
  input         clock, // @[:@3094.4]
  input         reset, // @[:@3095.4]
  input  [31:0] io_ibus_addr, // @[:@3096.4]
  output [31:0] io_ibus_inst, // @[:@3096.4]
  output        io_ibus_valid, // @[:@3096.4]
  input  [15:0] io_wbs_m2s_addr, // @[:@3096.4]
  input  [31:0] io_wbs_m2s_data, // @[:@3096.4]
  input         io_wbs_m2s_we, // @[:@3096.4]
  input  [3:0]  io_wbs_m2s_sel, // @[:@3096.4]
  input         io_wbs_m2s_stb, // @[:@3096.4]
  output        io_wbs_ack_o, // @[:@3096.4]
  output [31:0] io_wbs_data_o // @[:@3096.4]
);
  wire  imem_clock; // @[imem_interface.scala 40:20:@3098.4]
  wire [31:0] imem_io_imem_addr; // @[imem_interface.scala 40:20:@3098.4]
  wire [31:0] imem_io_imem_rdata; // @[imem_interface.scala 40:20:@3098.4]
  wire [31:0] imem_io_imem_wdata; // @[imem_interface.scala 40:20:@3098.4]
  wire  imem_io_wr_en; // @[imem_interface.scala 40:20:@3098.4]
  wire  bmem_clock; // @[imem_interface.scala 41:20:@3101.4]
  wire  bmem_reset; // @[imem_interface.scala 41:20:@3101.4]
  wire [31:0] bmem_io_bmem_addr; // @[imem_interface.scala 41:20:@3101.4]
  wire [31:0] bmem_io_bmem_rdata; // @[imem_interface.scala 41:20:@3101.4]
  wire [11:0] ibus_imem_addr; // @[imem_interface.scala 47:41:@3104.4]
  wire [11:0] wbs_imem_addr; // @[imem_interface.scala 49:44:@3106.4]
  reg  ack; // @[imem_interface.scala 54:31:@3107.4]
  reg [31:0] _RAND_0;
  reg [3:0] wb_select; // @[imem_interface.scala 55:27:@3108.4]
  reg [31:0] _RAND_1;
  wire  _T_45; // @[imem_interface.scala 57:24:@3109.4]
  wire  wb_rd_en; // @[imem_interface.scala 57:39:@3110.4]
  wire  wb_wr_en; // @[imem_interface.scala 58:38:@3111.4]
  wire [3:0] _T_46; // @[imem_interface.scala 63:46:@3112.4]
  wire  _T_48; // @[imem_interface.scala 63:84:@3113.4]
  wire  imem_wbs_addr_match; // @[imem_interface.scala 63:29:@3114.4]
  wire  _T_52; // @[imem_interface.scala 70:33:@3118.4]
  wire  imem_wbs_sel; // @[imem_interface.scala 70:46:@3119.4]
  reg  imem_ibus_valid; // @[imem_interface.scala 71:32:@3121.4]
  reg [31:0] _RAND_2;
  wire  _T_57; // @[imem_interface.scala 72:22:@3122.4]
  wire [11:0] imem_addr; // @[imem_interface.scala 80:27:@3128.4]
  wire [31:0] rd_imem_inst; // @[imem_interface.scala 92:23:@3133.4]
  wire [31:0] rd_imem_const; // @[imem_interface.scala 92:23:@3133.4]
  wire  _GEN_2; // @[imem_interface.scala 98:20:@3139.4]
  wire  _T_64; // @[imem_interface.scala 106:18:@3145.4]
  wire [7:0] _T_65; // @[imem_interface.scala 107:33:@3147.6]
  wire  _T_66; // @[imem_interface.scala 108:24:@3151.6]
  wire [7:0] _T_67; // @[imem_interface.scala 109:33:@3153.8]
  wire  _T_68; // @[imem_interface.scala 110:24:@3157.8]
  wire [7:0] _T_69; // @[imem_interface.scala 111:33:@3159.10]
  wire  _T_70; // @[imem_interface.scala 112:24:@3163.10]
  wire [7:0] _T_71; // @[imem_interface.scala 113:33:@3165.12]
  wire  _T_72; // @[imem_interface.scala 114:24:@3169.12]
  wire [15:0] _T_73; // @[imem_interface.scala 115:33:@3171.14]
  wire  _T_74; // @[imem_interface.scala 116:24:@3175.14]
  wire [15:0] _T_75; // @[imem_interface.scala 117:33:@3177.16]
  wire [31:0] _GEN_3; // @[imem_interface.scala 116:54:@3176.14]
  wire [31:0] _GEN_4; // @[imem_interface.scala 114:52:@3170.12]
  wire [31:0] _GEN_5; // @[imem_interface.scala 112:52:@3164.10]
  wire [31:0] _GEN_6; // @[imem_interface.scala 110:52:@3158.8]
  wire [31:0] _GEN_7; // @[imem_interface.scala 108:52:@3152.6]
  reg  bmem_ibus_sel; // @[imem_interface.scala 127:31:@3186.4]
  reg [31:0] _RAND_3;
  wire [3:0] _T_79; // @[imem_interface.scala 128:34:@3187.4]
  wire  _T_81; // @[imem_interface.scala 128:66:@3188.4]
  IMem imem ( // @[imem_interface.scala 40:20:@3098.4]
    .clock(imem_clock),
    .io_imem_addr(imem_io_imem_addr),
    .io_imem_rdata(imem_io_imem_rdata),
    .io_imem_wdata(imem_io_imem_wdata),
    .io_wr_en(imem_io_wr_en)
  );
  BMem bmem ( // @[imem_interface.scala 41:20:@3101.4]
    .clock(bmem_clock),
    .reset(bmem_reset),
    .io_bmem_addr(bmem_io_bmem_addr),
    .io_bmem_rdata(bmem_io_bmem_rdata)
  );
  assign ibus_imem_addr = io_ibus_addr[11:0]; // @[imem_interface.scala 47:41:@3104.4]
  assign wbs_imem_addr = io_wbs_m2s_addr[11:0]; // @[imem_interface.scala 49:44:@3106.4]
  assign _T_45 = io_wbs_m2s_we == 1'h0; // @[imem_interface.scala 57:24:@3109.4]
  assign wb_rd_en = _T_45 & io_wbs_m2s_stb; // @[imem_interface.scala 57:39:@3110.4]
  assign wb_wr_en = io_wbs_m2s_we & io_wbs_m2s_stb; // @[imem_interface.scala 58:38:@3111.4]
  assign _T_46 = io_wbs_m2s_addr[15:12]; // @[imem_interface.scala 63:46:@3112.4]
  assign _T_48 = _T_46 != 4'h0; // @[imem_interface.scala 63:84:@3113.4]
  assign imem_wbs_addr_match = _T_48 == 1'h0; // @[imem_interface.scala 63:29:@3114.4]
  assign _T_52 = wb_rd_en | wb_wr_en; // @[imem_interface.scala 70:33:@3118.4]
  assign imem_wbs_sel = _T_52 & imem_wbs_addr_match; // @[imem_interface.scala 70:46:@3119.4]
  assign _T_57 = imem_wbs_sel == 1'h0; // @[imem_interface.scala 72:22:@3122.4]
  assign imem_addr = imem_wbs_sel ? wbs_imem_addr : ibus_imem_addr; // @[imem_interface.scala 80:27:@3128.4]
  assign rd_imem_inst = imem_ibus_valid ? imem_io_imem_rdata : 32'h0; // @[imem_interface.scala 92:23:@3133.4]
  assign rd_imem_const = imem_ibus_valid ? 32'h0 : imem_io_imem_rdata; // @[imem_interface.scala 92:23:@3133.4]
  assign _GEN_2 = imem_wbs_sel ? io_wbs_m2s_stb : ack; // @[imem_interface.scala 98:20:@3139.4]
  assign _T_64 = wb_select == 4'h1; // @[imem_interface.scala 106:18:@3145.4]
  assign _T_65 = rd_imem_const[7:0]; // @[imem_interface.scala 107:33:@3147.6]
  assign _T_66 = wb_select == 4'h2; // @[imem_interface.scala 108:24:@3151.6]
  assign _T_67 = rd_imem_const[15:8]; // @[imem_interface.scala 109:33:@3153.8]
  assign _T_68 = wb_select == 4'h4; // @[imem_interface.scala 110:24:@3157.8]
  assign _T_69 = rd_imem_const[23:16]; // @[imem_interface.scala 111:33:@3159.10]
  assign _T_70 = wb_select == 4'h8; // @[imem_interface.scala 112:24:@3163.10]
  assign _T_71 = rd_imem_const[31:24]; // @[imem_interface.scala 113:33:@3165.12]
  assign _T_72 = wb_select == 4'h3; // @[imem_interface.scala 114:24:@3169.12]
  assign _T_73 = rd_imem_const[15:0]; // @[imem_interface.scala 115:33:@3171.14]
  assign _T_74 = wb_select == 4'hc; // @[imem_interface.scala 116:24:@3175.14]
  assign _T_75 = rd_imem_const[31:16]; // @[imem_interface.scala 117:33:@3177.16]
  assign _GEN_3 = _T_74 ? {{16'd0}, _T_75} : rd_imem_const; // @[imem_interface.scala 116:54:@3176.14]
  assign _GEN_4 = _T_72 ? {{16'd0}, _T_73} : _GEN_3; // @[imem_interface.scala 114:52:@3170.12]
  assign _GEN_5 = _T_70 ? {{24'd0}, _T_71} : _GEN_4; // @[imem_interface.scala 112:52:@3164.10]
  assign _GEN_6 = _T_68 ? {{24'd0}, _T_69} : _GEN_5; // @[imem_interface.scala 110:52:@3158.8]
  assign _GEN_7 = _T_66 ? {{24'd0}, _T_67} : _GEN_6; // @[imem_interface.scala 108:52:@3152.6]
  assign _T_79 = io_ibus_addr[15:12]; // @[imem_interface.scala 128:34:@3187.4]
  assign _T_81 = _T_79 == 4'h7; // @[imem_interface.scala 128:66:@3188.4]
  assign io_ibus_inst = bmem_ibus_sel ? bmem_io_bmem_rdata : rd_imem_inst; // @[imem_interface.scala 137:19:@3192.4]
  assign io_ibus_valid = bmem_ibus_sel ? 1'h1 : imem_ibus_valid; // @[imem_interface.scala 138:19:@3194.4]
  assign io_wbs_ack_o = ack; // @[imem_interface.scala 123:18:@3184.4]
  assign io_wbs_data_o = _T_64 ? {{24'd0}, _T_65} : _GEN_7; // @[imem_interface.scala 124:18:@3185.4]
  assign imem_clock = clock; // @[:@3099.4]
  assign imem_io_imem_addr = {{20'd0}, imem_addr}; // @[imem_interface.scala 81:21:@3129.4]
  assign imem_io_imem_wdata = io_wbs_m2s_data; // @[imem_interface.scala 87:22:@3130.4]
  assign imem_io_wr_en = imem_wbs_addr_match & wb_wr_en; // @[imem_interface.scala 88:17:@3131.4]
  assign bmem_clock = clock; // @[:@3102.4]
  assign bmem_reset = reset; // @[:@3103.4]
  assign bmem_io_bmem_addr = {{20'd0}, ibus_imem_addr}; // @[imem_interface.scala 130:21:@3190.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ack = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  wb_select = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  imem_ibus_valid = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  bmem_ibus_sel = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ack <= 1'h1;
    end else begin
      if (imem_wbs_sel) begin
        ack <= io_wbs_m2s_stb;
      end
    end
    wb_select <= io_wbs_m2s_sel;
    if (reset) begin
      imem_ibus_valid <= 1'h1;
    end else begin
      imem_ibus_valid <= _T_57;
    end
    if (reset) begin
      bmem_ibus_sel <= 1'h0;
    end else begin
      bmem_ibus_sel <= _T_81;
    end
  end
endmodule

module IMem( // @[:@1977.2]
  input         clock, // @[:@1978.4]
  input  [31:0] io_imem_addr, // @[:@1980.4]
  output [31:0] io_imem_rdata, // @[:@1980.4]
  input  [31:0] io_imem_wdata, // @[:@1980.4]
  input         io_wr_en // @[:@1980.4]
);
  reg [31:0] imem [0:4095]; // @[memory.scala 32:25:@1982.4]
  reg [31:0] _RAND_0;
  wire [31:0] imem__T_24_data; // @[memory.scala 32:25:@1982.4]
  wire [11:0] imem__T_24_addr; // @[memory.scala 32:25:@1982.4]
  wire [31:0] imem__T_20_data; // @[memory.scala 32:25:@1982.4]
  wire [11:0] imem__T_20_addr; // @[memory.scala 32:25:@1982.4]
  wire  imem__T_20_mask; // @[memory.scala 32:25:@1982.4]
  wire  imem__T_20_en; // @[memory.scala 32:25:@1982.4]
  wire [31:0] _T_18; // @[memory.scala 43:23:@1984.6]
  wire [11:0] _T_19; // @[memory.scala 43:9:@1985.6]
  wire  _GEN_3; // @[memory.scala 42:19:@1983.4]
  reg [11:0] imem__T_24_addr_pipe_0;
  reg [31:0] _RAND_1;
  assign imem__T_24_addr = imem__T_24_addr_pipe_0;
  assign imem__T_24_data = imem[imem__T_24_addr]; // @[memory.scala 32:25:@1982.4]
  assign imem__T_20_data = io_imem_wdata;
  assign imem__T_20_addr = _T_18[11:0];
  assign imem__T_20_mask = 1'h1;
  assign imem__T_20_en = io_wr_en;
  assign _T_18 = io_imem_addr / 32'h4; // @[memory.scala 43:23:@1984.6]
  assign _T_19 = _T_18[11:0]; // @[memory.scala 43:9:@1985.6]
  assign _GEN_3 = 1'h1; // @[memory.scala 42:19:@1983.4]
  assign io_imem_rdata = imem__T_24_data; // @[memory.scala 61:17:@1992.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4096; initvar = initvar+1)
    imem[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  imem__T_24_addr_pipe_0 = _RAND_1[11:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(imem__T_20_en & imem__T_20_mask) begin
      imem[imem__T_20_addr] <= imem__T_20_data; // @[memory.scala 32:25:@1982.4]
    end
    if (_GEN_3) begin
      imem__T_24_addr_pipe_0 <= _T_19;
    end
  end
endmodule

module BMem( // @[:@1994.2]
  input         clock, // @[:@1995.4]
  input         reset, // @[:@1996.4]
  input  [31:0] io_bmem_addr, // @[:@1997.4]
  output [31:0] io_bmem_rdata // @[:@1997.4]
);
  wire [9:0] _T_9; // @[BMEM.scala 24:26:@1999.4]
  wire [9:0] addr; // @[BMEM.scala 24:33:@2000.4]
  reg [31:0] bmem_data; // @[BMEM.scala 25:26:@2001.4]
  reg [31:0] _RAND_0;
  wire  _T_14; // @[Conditional.scala 37:30:@2002.4]
  wire  _T_17; // @[Conditional.scala 37:30:@2007.6]
  wire  _T_20; // @[Conditional.scala 37:30:@2012.8]
  wire  _T_23; // @[Conditional.scala 37:30:@2017.10]
  wire  _T_26; // @[Conditional.scala 37:30:@2022.12]
  wire  _T_29; // @[Conditional.scala 37:30:@2027.14]
  wire  _T_32; // @[Conditional.scala 37:30:@2032.16]
  wire  _T_35; // @[Conditional.scala 37:30:@2037.18]
  wire  _T_38; // @[Conditional.scala 37:30:@2042.20]
  wire  _T_41; // @[Conditional.scala 37:30:@2047.22]
  wire  _T_44; // @[Conditional.scala 37:30:@2052.24]
  wire  _T_47; // @[Conditional.scala 37:30:@2057.26]
  wire  _T_50; // @[Conditional.scala 37:30:@2062.28]
  wire  _T_53; // @[Conditional.scala 37:30:@2067.30]
  wire  _T_56; // @[Conditional.scala 37:30:@2072.32]
  wire  _T_59; // @[Conditional.scala 37:30:@2077.34]
  wire  _T_62; // @[Conditional.scala 37:30:@2082.36]
  wire  _T_65; // @[Conditional.scala 37:30:@2087.38]
  wire  _T_68; // @[Conditional.scala 37:30:@2092.40]
  wire  _T_71; // @[Conditional.scala 37:30:@2097.42]
  wire  _T_74; // @[Conditional.scala 37:30:@2102.44]
  wire  _T_77; // @[Conditional.scala 37:30:@2107.46]
  wire  _T_80; // @[Conditional.scala 37:30:@2112.48]
  wire  _T_83; // @[Conditional.scala 37:30:@2117.50]
  wire  _T_86; // @[Conditional.scala 37:30:@2122.52]
  wire  _T_89; // @[Conditional.scala 37:30:@2127.54]
  wire  _T_92; // @[Conditional.scala 37:30:@2132.56]
  wire  _T_95; // @[Conditional.scala 37:30:@2137.58]
  wire  _T_98; // @[Conditional.scala 37:30:@2142.60]
  wire  _T_101; // @[Conditional.scala 37:30:@2147.62]
  wire  _T_104; // @[Conditional.scala 37:30:@2152.64]
  wire  _T_107; // @[Conditional.scala 37:30:@2157.66]
  wire  _T_110; // @[Conditional.scala 37:30:@2162.68]
  wire  _T_113; // @[Conditional.scala 37:30:@2167.70]
  wire  _T_116; // @[Conditional.scala 37:30:@2172.72]
  wire  _T_119; // @[Conditional.scala 37:30:@2177.74]
  wire  _T_122; // @[Conditional.scala 37:30:@2182.76]
  wire  _T_125; // @[Conditional.scala 37:30:@2187.78]
  wire  _T_128; // @[Conditional.scala 37:30:@2192.80]
  wire  _T_131; // @[Conditional.scala 37:30:@2197.82]
  wire  _T_134; // @[Conditional.scala 37:30:@2202.84]
  wire  _T_137; // @[Conditional.scala 37:30:@2207.86]
  wire  _T_140; // @[Conditional.scala 37:30:@2212.88]
  wire  _T_143; // @[Conditional.scala 37:30:@2217.90]
  wire  _T_146; // @[Conditional.scala 37:30:@2222.92]
  wire  _T_149; // @[Conditional.scala 37:30:@2227.94]
  wire  _T_152; // @[Conditional.scala 37:30:@2232.96]
  wire  _T_155; // @[Conditional.scala 37:30:@2237.98]
  wire  _T_158; // @[Conditional.scala 37:30:@2242.100]
  wire  _T_161; // @[Conditional.scala 37:30:@2247.102]
  wire  _T_164; // @[Conditional.scala 37:30:@2252.104]
  wire  _T_167; // @[Conditional.scala 37:30:@2257.106]
  wire  _T_170; // @[Conditional.scala 37:30:@2262.108]
  wire  _T_173; // @[Conditional.scala 37:30:@2267.110]
  wire  _T_176; // @[Conditional.scala 37:30:@2272.112]
  wire  _T_179; // @[Conditional.scala 37:30:@2277.114]
  wire  _T_182; // @[Conditional.scala 37:30:@2282.116]
  wire  _T_185; // @[Conditional.scala 37:30:@2287.118]
  wire  _T_188; // @[Conditional.scala 37:30:@2292.120]
  wire  _T_191; // @[Conditional.scala 37:30:@2297.122]
  wire  _T_194; // @[Conditional.scala 37:30:@2302.124]
  wire  _T_197; // @[Conditional.scala 37:30:@2307.126]
  wire  _T_200; // @[Conditional.scala 37:30:@2312.128]
  wire  _T_203; // @[Conditional.scala 37:30:@2317.130]
  wire  _T_206; // @[Conditional.scala 37:30:@2322.132]
  wire  _T_209; // @[Conditional.scala 37:30:@2327.134]
  wire  _T_212; // @[Conditional.scala 37:30:@2332.136]
  wire  _T_215; // @[Conditional.scala 37:30:@2337.138]
  wire  _T_218; // @[Conditional.scala 37:30:@2342.140]
  wire  _T_221; // @[Conditional.scala 37:30:@2347.142]
  wire  _T_224; // @[Conditional.scala 37:30:@2352.144]
  wire  _T_227; // @[Conditional.scala 37:30:@2357.146]
  wire  _T_230; // @[Conditional.scala 37:30:@2362.148]
  wire  _T_233; // @[Conditional.scala 37:30:@2367.150]
  wire  _T_236; // @[Conditional.scala 37:30:@2372.152]
  wire  _T_239; // @[Conditional.scala 37:30:@2377.154]
  wire  _T_242; // @[Conditional.scala 37:30:@2382.156]
  wire  _T_245; // @[Conditional.scala 37:30:@2387.158]
  wire  _T_248; // @[Conditional.scala 37:30:@2392.160]
  wire  _T_251; // @[Conditional.scala 37:30:@2397.162]
  wire  _T_254; // @[Conditional.scala 37:30:@2402.164]
  wire  _T_257; // @[Conditional.scala 37:30:@2407.166]
  wire  _T_260; // @[Conditional.scala 37:30:@2412.168]
  wire  _T_263; // @[Conditional.scala 37:30:@2417.170]
  wire  _T_266; // @[Conditional.scala 37:30:@2422.172]
  wire  _T_269; // @[Conditional.scala 37:30:@2427.174]
  wire  _T_272; // @[Conditional.scala 37:30:@2432.176]
  wire  _T_275; // @[Conditional.scala 37:30:@2437.178]
  wire  _T_278; // @[Conditional.scala 37:30:@2442.180]
  wire  _T_281; // @[Conditional.scala 37:30:@2447.182]
  wire  _T_284; // @[Conditional.scala 37:30:@2452.184]
  wire  _T_287; // @[Conditional.scala 37:30:@2457.186]
  wire  _T_290; // @[Conditional.scala 37:30:@2462.188]
  wire  _T_293; // @[Conditional.scala 37:30:@2467.190]
  wire  _T_296; // @[Conditional.scala 37:30:@2472.192]
  wire  _T_299; // @[Conditional.scala 37:30:@2477.194]
  wire  _T_302; // @[Conditional.scala 37:30:@2482.196]
  wire  _T_305; // @[Conditional.scala 37:30:@2487.198]
  wire  _T_308; // @[Conditional.scala 37:30:@2492.200]
  wire  _T_311; // @[Conditional.scala 37:30:@2497.202]
  wire  _T_314; // @[Conditional.scala 37:30:@2502.204]
  wire  _T_317; // @[Conditional.scala 37:30:@2507.206]
  wire  _T_320; // @[Conditional.scala 37:30:@2512.208]
  wire  _T_323; // @[Conditional.scala 37:30:@2517.210]
  wire  _T_326; // @[Conditional.scala 37:30:@2522.212]
  wire  _T_329; // @[Conditional.scala 37:30:@2527.214]
  wire  _T_332; // @[Conditional.scala 37:30:@2532.216]
  wire  _T_335; // @[Conditional.scala 37:30:@2537.218]
  wire  _T_338; // @[Conditional.scala 37:30:@2542.220]
  wire  _T_341; // @[Conditional.scala 37:30:@2547.222]
  wire  _T_344; // @[Conditional.scala 37:30:@2552.224]
  wire  _T_347; // @[Conditional.scala 37:30:@2557.226]
  wire  _T_350; // @[Conditional.scala 37:30:@2562.228]
  wire  _T_353; // @[Conditional.scala 37:30:@2567.230]
  wire  _T_356; // @[Conditional.scala 37:30:@2572.232]
  wire  _T_359; // @[Conditional.scala 37:30:@2577.234]
  wire  _T_362; // @[Conditional.scala 37:30:@2582.236]
  wire  _T_365; // @[Conditional.scala 37:30:@2587.238]
  wire  _T_368; // @[Conditional.scala 37:30:@2592.240]
  wire  _T_371; // @[Conditional.scala 37:30:@2597.242]
  wire  _T_374; // @[Conditional.scala 37:30:@2602.244]
  wire  _T_377; // @[Conditional.scala 37:30:@2607.246]
  wire  _T_380; // @[Conditional.scala 37:30:@2612.248]
  wire  _T_383; // @[Conditional.scala 37:30:@2617.250]
  wire  _T_386; // @[Conditional.scala 37:30:@2622.252]
  wire  _T_389; // @[Conditional.scala 37:30:@2627.254]
  wire  _T_392; // @[Conditional.scala 37:30:@2632.256]
  wire  _T_395; // @[Conditional.scala 37:30:@2637.258]
  wire  _T_398; // @[Conditional.scala 37:30:@2642.260]
  wire  _T_401; // @[Conditional.scala 37:30:@2647.262]
  wire  _T_404; // @[Conditional.scala 37:30:@2652.264]
  wire  _T_407; // @[Conditional.scala 37:30:@2657.266]
  wire  _T_410; // @[Conditional.scala 37:30:@2662.268]
  wire  _T_413; // @[Conditional.scala 37:30:@2667.270]
  wire  _T_416; // @[Conditional.scala 37:30:@2672.272]
  wire  _T_419; // @[Conditional.scala 37:30:@2677.274]
  wire  _T_422; // @[Conditional.scala 37:30:@2682.276]
  wire  _T_425; // @[Conditional.scala 37:30:@2687.278]
  wire  _T_428; // @[Conditional.scala 37:30:@2692.280]
  wire  _T_431; // @[Conditional.scala 37:30:@2697.282]
  wire  _T_434; // @[Conditional.scala 37:30:@2702.284]
  wire  _T_437; // @[Conditional.scala 37:30:@2707.286]
  wire  _T_440; // @[Conditional.scala 37:30:@2712.288]
  wire  _T_443; // @[Conditional.scala 37:30:@2717.290]
  wire  _T_446; // @[Conditional.scala 37:30:@2722.292]
  wire  _T_449; // @[Conditional.scala 37:30:@2727.294]
  wire  _T_452; // @[Conditional.scala 37:30:@2732.296]
  wire  _T_455; // @[Conditional.scala 37:30:@2737.298]
  wire  _T_458; // @[Conditional.scala 37:30:@2742.300]
  wire  _T_461; // @[Conditional.scala 37:30:@2747.302]
  wire  _T_464; // @[Conditional.scala 37:30:@2752.304]
  wire  _T_467; // @[Conditional.scala 37:30:@2757.306]
  wire  _T_470; // @[Conditional.scala 37:30:@2762.308]
  wire  _T_473; // @[Conditional.scala 37:30:@2767.310]
  wire  _T_476; // @[Conditional.scala 37:30:@2772.312]
  wire  _T_479; // @[Conditional.scala 37:30:@2777.314]
  wire  _T_482; // @[Conditional.scala 37:30:@2782.316]
  wire  _T_485; // @[Conditional.scala 37:30:@2787.318]
  wire  _T_488; // @[Conditional.scala 37:30:@2792.320]
  wire  _T_491; // @[Conditional.scala 37:30:@2797.322]
  wire  _T_494; // @[Conditional.scala 37:30:@2802.324]
  wire  _T_497; // @[Conditional.scala 37:30:@2807.326]
  wire  _T_500; // @[Conditional.scala 37:30:@2812.328]
  wire  _T_503; // @[Conditional.scala 37:30:@2817.330]
  wire  _T_506; // @[Conditional.scala 37:30:@2822.332]
  wire  _T_509; // @[Conditional.scala 37:30:@2827.334]
  wire  _T_512; // @[Conditional.scala 37:30:@2832.336]
  wire  _T_515; // @[Conditional.scala 37:30:@2837.338]
  wire  _T_518; // @[Conditional.scala 37:30:@2842.340]
  wire  _T_521; // @[Conditional.scala 37:30:@2847.342]
  wire  _T_524; // @[Conditional.scala 37:30:@2852.344]
  wire  _T_527; // @[Conditional.scala 37:30:@2857.346]
  wire  _T_530; // @[Conditional.scala 37:30:@2862.348]
  wire  _T_533; // @[Conditional.scala 37:30:@2867.350]
  wire  _T_536; // @[Conditional.scala 37:30:@2872.352]
  wire  _T_539; // @[Conditional.scala 37:30:@2877.354]
  wire  _T_542; // @[Conditional.scala 37:30:@2882.356]
  wire  _T_545; // @[Conditional.scala 37:30:@2887.358]
  wire  _T_548; // @[Conditional.scala 37:30:@2892.360]
  wire  _T_551; // @[Conditional.scala 37:30:@2897.362]
  wire  _T_554; // @[Conditional.scala 37:30:@2902.364]
  wire  _T_557; // @[Conditional.scala 37:30:@2907.366]
  wire  _T_560; // @[Conditional.scala 37:30:@2912.368]
  wire  _T_563; // @[Conditional.scala 37:30:@2917.370]
  wire  _T_566; // @[Conditional.scala 37:30:@2922.372]
  wire  _T_569; // @[Conditional.scala 37:30:@2927.374]
  wire  _T_572; // @[Conditional.scala 37:30:@2932.376]
  wire  _T_575; // @[Conditional.scala 37:30:@2937.378]
  wire  _T_578; // @[Conditional.scala 37:30:@2942.380]
  wire  _T_581; // @[Conditional.scala 37:30:@2947.382]
  wire  _T_584; // @[Conditional.scala 37:30:@2952.384]
  wire  _T_587; // @[Conditional.scala 37:30:@2957.386]
  wire  _T_590; // @[Conditional.scala 37:30:@2962.388]
  wire  _T_593; // @[Conditional.scala 37:30:@2967.390]
  wire  _T_596; // @[Conditional.scala 37:30:@2972.392]
  wire  _T_599; // @[Conditional.scala 37:30:@2977.394]
  wire  _T_602; // @[Conditional.scala 37:30:@2982.396]
  wire  _T_605; // @[Conditional.scala 37:30:@2987.398]
  wire  _T_608; // @[Conditional.scala 37:30:@2992.400]
  wire  _T_611; // @[Conditional.scala 37:30:@2997.402]
  wire  _T_614; // @[Conditional.scala 37:30:@3002.404]
  wire  _T_617; // @[Conditional.scala 37:30:@3007.406]
  wire  _T_620; // @[Conditional.scala 37:30:@3012.408]
  wire  _T_623; // @[Conditional.scala 37:30:@3017.410]
  wire  _T_626; // @[Conditional.scala 37:30:@3022.412]
  wire  _T_629; // @[Conditional.scala 37:30:@3027.414]
  wire  _T_632; // @[Conditional.scala 37:30:@3032.416]
  wire  _T_635; // @[Conditional.scala 37:30:@3037.418]
  wire  _T_638; // @[Conditional.scala 37:30:@3042.420]
  wire  _T_641; // @[Conditional.scala 37:30:@3047.422]
  wire  _T_644; // @[Conditional.scala 37:30:@3052.424]
  wire  _T_647; // @[Conditional.scala 37:30:@3057.426]
  wire  _T_650; // @[Conditional.scala 37:30:@3062.428]
  wire  _T_653; // @[Conditional.scala 37:30:@3067.430]
  wire  _T_656; // @[Conditional.scala 37:30:@3072.432]
  wire  _T_659; // @[Conditional.scala 37:30:@3077.434]
  wire  _T_662; // @[Conditional.scala 37:30:@3082.436]
  wire  _T_665; // @[Conditional.scala 37:30:@3087.438]
  wire [31:0] _GEN_0; // @[Conditional.scala 39:67:@3088.438]
  wire [31:0] _GEN_1; // @[Conditional.scala 39:67:@3083.436]
  wire [31:0] _GEN_2; // @[Conditional.scala 39:67:@3078.434]
  wire [31:0] _GEN_3; // @[Conditional.scala 39:67:@3073.432]
  wire [31:0] _GEN_4; // @[Conditional.scala 39:67:@3068.430]
  wire [31:0] _GEN_5; // @[Conditional.scala 39:67:@3063.428]
  wire [31:0] _GEN_6; // @[Conditional.scala 39:67:@3058.426]
  wire [31:0] _GEN_7; // @[Conditional.scala 39:67:@3053.424]
  wire [31:0] _GEN_8; // @[Conditional.scala 39:67:@3048.422]
  wire [31:0] _GEN_9; // @[Conditional.scala 39:67:@3043.420]
  wire [31:0] _GEN_10; // @[Conditional.scala 39:67:@3038.418]
  wire [31:0] _GEN_11; // @[Conditional.scala 39:67:@3033.416]
  wire [31:0] _GEN_12; // @[Conditional.scala 39:67:@3028.414]
  wire [31:0] _GEN_13; // @[Conditional.scala 39:67:@3023.412]
  wire [31:0] _GEN_14; // @[Conditional.scala 39:67:@3018.410]
  wire [31:0] _GEN_15; // @[Conditional.scala 39:67:@3013.408]
  wire [31:0] _GEN_16; // @[Conditional.scala 39:67:@3008.406]
  wire [31:0] _GEN_17; // @[Conditional.scala 39:67:@3003.404]
  wire [31:0] _GEN_18; // @[Conditional.scala 39:67:@2998.402]
  wire [31:0] _GEN_19; // @[Conditional.scala 39:67:@2993.400]
  wire [31:0] _GEN_20; // @[Conditional.scala 39:67:@2988.398]
  wire [31:0] _GEN_21; // @[Conditional.scala 39:67:@2983.396]
  wire [31:0] _GEN_22; // @[Conditional.scala 39:67:@2978.394]
  wire [31:0] _GEN_23; // @[Conditional.scala 39:67:@2973.392]
  wire [31:0] _GEN_24; // @[Conditional.scala 39:67:@2968.390]
  wire [31:0] _GEN_25; // @[Conditional.scala 39:67:@2963.388]
  wire [31:0] _GEN_26; // @[Conditional.scala 39:67:@2958.386]
  wire [31:0] _GEN_27; // @[Conditional.scala 39:67:@2953.384]
  wire [31:0] _GEN_28; // @[Conditional.scala 39:67:@2948.382]
  wire [31:0] _GEN_29; // @[Conditional.scala 39:67:@2943.380]
  wire [31:0] _GEN_30; // @[Conditional.scala 39:67:@2938.378]
  wire [31:0] _GEN_31; // @[Conditional.scala 39:67:@2933.376]
  wire [31:0] _GEN_32; // @[Conditional.scala 39:67:@2928.374]
  wire [31:0] _GEN_33; // @[Conditional.scala 39:67:@2923.372]
  wire [31:0] _GEN_34; // @[Conditional.scala 39:67:@2918.370]
  wire [31:0] _GEN_35; // @[Conditional.scala 39:67:@2913.368]
  wire [31:0] _GEN_36; // @[Conditional.scala 39:67:@2908.366]
  wire [31:0] _GEN_37; // @[Conditional.scala 39:67:@2903.364]
  wire [31:0] _GEN_38; // @[Conditional.scala 39:67:@2898.362]
  wire [31:0] _GEN_39; // @[Conditional.scala 39:67:@2893.360]
  wire [31:0] _GEN_40; // @[Conditional.scala 39:67:@2888.358]
  wire [31:0] _GEN_41; // @[Conditional.scala 39:67:@2883.356]
  wire [31:0] _GEN_42; // @[Conditional.scala 39:67:@2878.354]
  wire [31:0] _GEN_43; // @[Conditional.scala 39:67:@2873.352]
  wire [31:0] _GEN_44; // @[Conditional.scala 39:67:@2868.350]
  wire [31:0] _GEN_45; // @[Conditional.scala 39:67:@2863.348]
  wire [31:0] _GEN_46; // @[Conditional.scala 39:67:@2858.346]
  wire [31:0] _GEN_47; // @[Conditional.scala 39:67:@2853.344]
  wire [31:0] _GEN_48; // @[Conditional.scala 39:67:@2848.342]
  wire [31:0] _GEN_49; // @[Conditional.scala 39:67:@2843.340]
  wire [31:0] _GEN_50; // @[Conditional.scala 39:67:@2838.338]
  wire [31:0] _GEN_51; // @[Conditional.scala 39:67:@2833.336]
  wire [31:0] _GEN_52; // @[Conditional.scala 39:67:@2828.334]
  wire [31:0] _GEN_53; // @[Conditional.scala 39:67:@2823.332]
  wire [31:0] _GEN_54; // @[Conditional.scala 39:67:@2818.330]
  wire [31:0] _GEN_55; // @[Conditional.scala 39:67:@2813.328]
  wire [31:0] _GEN_56; // @[Conditional.scala 39:67:@2808.326]
  wire [31:0] _GEN_57; // @[Conditional.scala 39:67:@2803.324]
  wire [31:0] _GEN_58; // @[Conditional.scala 39:67:@2798.322]
  wire [31:0] _GEN_59; // @[Conditional.scala 39:67:@2793.320]
  wire [31:0] _GEN_60; // @[Conditional.scala 39:67:@2788.318]
  wire [31:0] _GEN_61; // @[Conditional.scala 39:67:@2783.316]
  wire [31:0] _GEN_62; // @[Conditional.scala 39:67:@2778.314]
  wire [31:0] _GEN_63; // @[Conditional.scala 39:67:@2773.312]
  wire [31:0] _GEN_64; // @[Conditional.scala 39:67:@2768.310]
  wire [31:0] _GEN_65; // @[Conditional.scala 39:67:@2763.308]
  wire [31:0] _GEN_66; // @[Conditional.scala 39:67:@2758.306]
  wire [31:0] _GEN_67; // @[Conditional.scala 39:67:@2753.304]
  wire [31:0] _GEN_68; // @[Conditional.scala 39:67:@2748.302]
  wire [31:0] _GEN_69; // @[Conditional.scala 39:67:@2743.300]
  wire [31:0] _GEN_70; // @[Conditional.scala 39:67:@2738.298]
  wire [31:0] _GEN_71; // @[Conditional.scala 39:67:@2733.296]
  wire [31:0] _GEN_72; // @[Conditional.scala 39:67:@2728.294]
  wire [31:0] _GEN_73; // @[Conditional.scala 39:67:@2723.292]
  wire [31:0] _GEN_74; // @[Conditional.scala 39:67:@2718.290]
  wire [31:0] _GEN_75; // @[Conditional.scala 39:67:@2713.288]
  wire [31:0] _GEN_76; // @[Conditional.scala 39:67:@2708.286]
  wire [31:0] _GEN_77; // @[Conditional.scala 39:67:@2703.284]
  wire [31:0] _GEN_78; // @[Conditional.scala 39:67:@2698.282]
  wire [31:0] _GEN_79; // @[Conditional.scala 39:67:@2693.280]
  wire [31:0] _GEN_80; // @[Conditional.scala 39:67:@2688.278]
  wire [31:0] _GEN_81; // @[Conditional.scala 39:67:@2683.276]
  wire [31:0] _GEN_82; // @[Conditional.scala 39:67:@2678.274]
  wire [31:0] _GEN_83; // @[Conditional.scala 39:67:@2673.272]
  wire [31:0] _GEN_84; // @[Conditional.scala 39:67:@2668.270]
  wire [31:0] _GEN_85; // @[Conditional.scala 39:67:@2663.268]
  wire [31:0] _GEN_86; // @[Conditional.scala 39:67:@2658.266]
  wire [31:0] _GEN_87; // @[Conditional.scala 39:67:@2653.264]
  wire [31:0] _GEN_88; // @[Conditional.scala 39:67:@2648.262]
  wire [31:0] _GEN_89; // @[Conditional.scala 39:67:@2643.260]
  wire [31:0] _GEN_90; // @[Conditional.scala 39:67:@2638.258]
  wire [31:0] _GEN_91; // @[Conditional.scala 39:67:@2633.256]
  wire [31:0] _GEN_92; // @[Conditional.scala 39:67:@2628.254]
  wire [31:0] _GEN_93; // @[Conditional.scala 39:67:@2623.252]
  wire [31:0] _GEN_94; // @[Conditional.scala 39:67:@2618.250]
  wire [31:0] _GEN_95; // @[Conditional.scala 39:67:@2613.248]
  wire [31:0] _GEN_96; // @[Conditional.scala 39:67:@2608.246]
  wire [31:0] _GEN_97; // @[Conditional.scala 39:67:@2603.244]
  wire [31:0] _GEN_98; // @[Conditional.scala 39:67:@2598.242]
  wire [31:0] _GEN_99; // @[Conditional.scala 39:67:@2593.240]
  wire [31:0] _GEN_100; // @[Conditional.scala 39:67:@2588.238]
  wire [31:0] _GEN_101; // @[Conditional.scala 39:67:@2583.236]
  wire [31:0] _GEN_102; // @[Conditional.scala 39:67:@2578.234]
  wire [31:0] _GEN_103; // @[Conditional.scala 39:67:@2573.232]
  wire [31:0] _GEN_104; // @[Conditional.scala 39:67:@2568.230]
  wire [31:0] _GEN_105; // @[Conditional.scala 39:67:@2563.228]
  wire [31:0] _GEN_106; // @[Conditional.scala 39:67:@2558.226]
  wire [31:0] _GEN_107; // @[Conditional.scala 39:67:@2553.224]
  wire [31:0] _GEN_108; // @[Conditional.scala 39:67:@2548.222]
  wire [31:0] _GEN_109; // @[Conditional.scala 39:67:@2543.220]
  wire [31:0] _GEN_110; // @[Conditional.scala 39:67:@2538.218]
  wire [31:0] _GEN_111; // @[Conditional.scala 39:67:@2533.216]
  wire [31:0] _GEN_112; // @[Conditional.scala 39:67:@2528.214]
  wire [31:0] _GEN_113; // @[Conditional.scala 39:67:@2523.212]
  wire [31:0] _GEN_114; // @[Conditional.scala 39:67:@2518.210]
  wire [31:0] _GEN_115; // @[Conditional.scala 39:67:@2513.208]
  wire [31:0] _GEN_116; // @[Conditional.scala 39:67:@2508.206]
  wire [31:0] _GEN_117; // @[Conditional.scala 39:67:@2503.204]
  wire [31:0] _GEN_118; // @[Conditional.scala 39:67:@2498.202]
  wire [31:0] _GEN_119; // @[Conditional.scala 39:67:@2493.200]
  wire [31:0] _GEN_120; // @[Conditional.scala 39:67:@2488.198]
  wire [31:0] _GEN_121; // @[Conditional.scala 39:67:@2483.196]
  wire [31:0] _GEN_122; // @[Conditional.scala 39:67:@2478.194]
  wire [31:0] _GEN_123; // @[Conditional.scala 39:67:@2473.192]
  wire [31:0] _GEN_124; // @[Conditional.scala 39:67:@2468.190]
  wire [31:0] _GEN_125; // @[Conditional.scala 39:67:@2463.188]
  wire [31:0] _GEN_126; // @[Conditional.scala 39:67:@2458.186]
  wire [31:0] _GEN_127; // @[Conditional.scala 39:67:@2453.184]
  wire [31:0] _GEN_128; // @[Conditional.scala 39:67:@2448.182]
  wire [31:0] _GEN_129; // @[Conditional.scala 39:67:@2443.180]
  wire [31:0] _GEN_130; // @[Conditional.scala 39:67:@2438.178]
  wire [31:0] _GEN_131; // @[Conditional.scala 39:67:@2433.176]
  wire [31:0] _GEN_132; // @[Conditional.scala 39:67:@2428.174]
  wire [31:0] _GEN_133; // @[Conditional.scala 39:67:@2423.172]
  wire [31:0] _GEN_134; // @[Conditional.scala 39:67:@2418.170]
  wire [31:0] _GEN_135; // @[Conditional.scala 39:67:@2413.168]
  wire [31:0] _GEN_136; // @[Conditional.scala 39:67:@2408.166]
  wire [31:0] _GEN_137; // @[Conditional.scala 39:67:@2403.164]
  wire [31:0] _GEN_138; // @[Conditional.scala 39:67:@2398.162]
  wire [31:0] _GEN_139; // @[Conditional.scala 39:67:@2393.160]
  wire [31:0] _GEN_140; // @[Conditional.scala 39:67:@2388.158]
  wire [31:0] _GEN_141; // @[Conditional.scala 39:67:@2383.156]
  wire [31:0] _GEN_142; // @[Conditional.scala 39:67:@2378.154]
  wire [31:0] _GEN_143; // @[Conditional.scala 39:67:@2373.152]
  wire [31:0] _GEN_144; // @[Conditional.scala 39:67:@2368.150]
  wire [31:0] _GEN_145; // @[Conditional.scala 39:67:@2363.148]
  wire [31:0] _GEN_146; // @[Conditional.scala 39:67:@2358.146]
  wire [31:0] _GEN_147; // @[Conditional.scala 39:67:@2353.144]
  wire [31:0] _GEN_148; // @[Conditional.scala 39:67:@2348.142]
  wire [31:0] _GEN_149; // @[Conditional.scala 39:67:@2343.140]
  wire [31:0] _GEN_150; // @[Conditional.scala 39:67:@2338.138]
  wire [31:0] _GEN_151; // @[Conditional.scala 39:67:@2333.136]
  wire [31:0] _GEN_152; // @[Conditional.scala 39:67:@2328.134]
  wire [31:0] _GEN_153; // @[Conditional.scala 39:67:@2323.132]
  wire [31:0] _GEN_154; // @[Conditional.scala 39:67:@2318.130]
  wire [31:0] _GEN_155; // @[Conditional.scala 39:67:@2313.128]
  wire [31:0] _GEN_156; // @[Conditional.scala 39:67:@2308.126]
  wire [31:0] _GEN_157; // @[Conditional.scala 39:67:@2303.124]
  wire [31:0] _GEN_158; // @[Conditional.scala 39:67:@2298.122]
  wire [31:0] _GEN_159; // @[Conditional.scala 39:67:@2293.120]
  wire [31:0] _GEN_160; // @[Conditional.scala 39:67:@2288.118]
  wire [31:0] _GEN_161; // @[Conditional.scala 39:67:@2283.116]
  wire [31:0] _GEN_162; // @[Conditional.scala 39:67:@2278.114]
  wire [31:0] _GEN_163; // @[Conditional.scala 39:67:@2273.112]
  wire [31:0] _GEN_164; // @[Conditional.scala 39:67:@2268.110]
  wire [31:0] _GEN_165; // @[Conditional.scala 39:67:@2263.108]
  wire [31:0] _GEN_166; // @[Conditional.scala 39:67:@2258.106]
  wire [31:0] _GEN_167; // @[Conditional.scala 39:67:@2253.104]
  wire [31:0] _GEN_168; // @[Conditional.scala 39:67:@2248.102]
  wire [31:0] _GEN_169; // @[Conditional.scala 39:67:@2243.100]
  wire [31:0] _GEN_170; // @[Conditional.scala 39:67:@2238.98]
  wire [31:0] _GEN_171; // @[Conditional.scala 39:67:@2233.96]
  wire [31:0] _GEN_172; // @[Conditional.scala 39:67:@2228.94]
  wire [31:0] _GEN_173; // @[Conditional.scala 39:67:@2223.92]
  wire [31:0] _GEN_174; // @[Conditional.scala 39:67:@2218.90]
  wire [31:0] _GEN_175; // @[Conditional.scala 39:67:@2213.88]
  wire [31:0] _GEN_176; // @[Conditional.scala 39:67:@2208.86]
  wire [31:0] _GEN_177; // @[Conditional.scala 39:67:@2203.84]
  wire [31:0] _GEN_178; // @[Conditional.scala 39:67:@2198.82]
  wire [31:0] _GEN_179; // @[Conditional.scala 39:67:@2193.80]
  wire [31:0] _GEN_180; // @[Conditional.scala 39:67:@2188.78]
  wire [31:0] _GEN_181; // @[Conditional.scala 39:67:@2183.76]
  wire [31:0] _GEN_182; // @[Conditional.scala 39:67:@2178.74]
  wire [31:0] _GEN_183; // @[Conditional.scala 39:67:@2173.72]
  wire [31:0] _GEN_184; // @[Conditional.scala 39:67:@2168.70]
  wire [31:0] _GEN_185; // @[Conditional.scala 39:67:@2163.68]
  wire [31:0] _GEN_186; // @[Conditional.scala 39:67:@2158.66]
  wire [31:0] _GEN_187; // @[Conditional.scala 39:67:@2153.64]
  wire [31:0] _GEN_188; // @[Conditional.scala 39:67:@2148.62]
  wire [31:0] _GEN_189; // @[Conditional.scala 39:67:@2143.60]
  wire [31:0] _GEN_190; // @[Conditional.scala 39:67:@2138.58]
  wire [31:0] _GEN_191; // @[Conditional.scala 39:67:@2133.56]
  wire [31:0] _GEN_192; // @[Conditional.scala 39:67:@2128.54]
  wire [31:0] _GEN_193; // @[Conditional.scala 39:67:@2123.52]
  wire [31:0] _GEN_194; // @[Conditional.scala 39:67:@2118.50]
  wire [31:0] _GEN_195; // @[Conditional.scala 39:67:@2113.48]
  wire [31:0] _GEN_196; // @[Conditional.scala 39:67:@2108.46]
  wire [31:0] _GEN_197; // @[Conditional.scala 39:67:@2103.44]
  wire [31:0] _GEN_198; // @[Conditional.scala 39:67:@2098.42]
  wire [31:0] _GEN_199; // @[Conditional.scala 39:67:@2093.40]
  wire [31:0] _GEN_200; // @[Conditional.scala 39:67:@2088.38]
  wire [31:0] _GEN_201; // @[Conditional.scala 39:67:@2083.36]
  wire [31:0] _GEN_202; // @[Conditional.scala 39:67:@2078.34]
  wire [31:0] _GEN_203; // @[Conditional.scala 39:67:@2073.32]
  wire [31:0] _GEN_204; // @[Conditional.scala 39:67:@2068.30]
  wire [31:0] _GEN_205; // @[Conditional.scala 39:67:@2063.28]
  wire [31:0] _GEN_206; // @[Conditional.scala 39:67:@2058.26]
  wire [31:0] _GEN_207; // @[Conditional.scala 39:67:@2053.24]
  wire [31:0] _GEN_208; // @[Conditional.scala 39:67:@2048.22]
  wire [31:0] _GEN_209; // @[Conditional.scala 39:67:@2043.20]
  wire [31:0] _GEN_210; // @[Conditional.scala 39:67:@2038.18]
  wire [31:0] _GEN_211; // @[Conditional.scala 39:67:@2033.16]
  wire [31:0] _GEN_212; // @[Conditional.scala 39:67:@2028.14]
  wire [31:0] _GEN_213; // @[Conditional.scala 39:67:@2023.12]
  wire [31:0] _GEN_214; // @[Conditional.scala 39:67:@2018.10]
  wire [31:0] _GEN_215; // @[Conditional.scala 39:67:@2013.8]
  wire [31:0] _GEN_216; // @[Conditional.scala 39:67:@2008.6]
  wire [31:0] _GEN_217; // @[Conditional.scala 40:58:@2003.4]
  assign _T_9 = io_bmem_addr[9:0]; // @[BMEM.scala 24:26:@1999.4]
  assign addr = _T_9 / 10'h4; // @[BMEM.scala 24:33:@2000.4]
  assign _T_14 = 10'h0 == addr; // @[Conditional.scala 37:30:@2002.4]
  assign _T_17 = 10'h1 == addr; // @[Conditional.scala 37:30:@2007.6]
  assign _T_20 = 10'h2 == addr; // @[Conditional.scala 37:30:@2012.8]
  assign _T_23 = 10'h3 == addr; // @[Conditional.scala 37:30:@2017.10]
  assign _T_26 = 10'h4 == addr; // @[Conditional.scala 37:30:@2022.12]
  assign _T_29 = 10'h5 == addr; // @[Conditional.scala 37:30:@2027.14]
  assign _T_32 = 10'h6 == addr; // @[Conditional.scala 37:30:@2032.16]
  assign _T_35 = 10'h7 == addr; // @[Conditional.scala 37:30:@2037.18]
  assign _T_38 = 10'h8 == addr; // @[Conditional.scala 37:30:@2042.20]
  assign _T_41 = 10'h9 == addr; // @[Conditional.scala 37:30:@2047.22]
  assign _T_44 = 10'ha == addr; // @[Conditional.scala 37:30:@2052.24]
  assign _T_47 = 10'hb == addr; // @[Conditional.scala 37:30:@2057.26]
  assign _T_50 = 10'hc == addr; // @[Conditional.scala 37:30:@2062.28]
  assign _T_53 = 10'hd == addr; // @[Conditional.scala 37:30:@2067.30]
  assign _T_56 = 10'he == addr; // @[Conditional.scala 37:30:@2072.32]
  assign _T_59 = 10'hf == addr; // @[Conditional.scala 37:30:@2077.34]
  assign _T_62 = 10'h10 == addr; // @[Conditional.scala 37:30:@2082.36]
  assign _T_65 = 10'h11 == addr; // @[Conditional.scala 37:30:@2087.38]
  assign _T_68 = 10'h12 == addr; // @[Conditional.scala 37:30:@2092.40]
  assign _T_71 = 10'h13 == addr; // @[Conditional.scala 37:30:@2097.42]
  assign _T_74 = 10'h14 == addr; // @[Conditional.scala 37:30:@2102.44]
  assign _T_77 = 10'h15 == addr; // @[Conditional.scala 37:30:@2107.46]
  assign _T_80 = 10'h16 == addr; // @[Conditional.scala 37:30:@2112.48]
  assign _T_83 = 10'h17 == addr; // @[Conditional.scala 37:30:@2117.50]
  assign _T_86 = 10'h18 == addr; // @[Conditional.scala 37:30:@2122.52]
  assign _T_89 = 10'h19 == addr; // @[Conditional.scala 37:30:@2127.54]
  assign _T_92 = 10'h1a == addr; // @[Conditional.scala 37:30:@2132.56]
  assign _T_95 = 10'h1b == addr; // @[Conditional.scala 37:30:@2137.58]
  assign _T_98 = 10'h1c == addr; // @[Conditional.scala 37:30:@2142.60]
  assign _T_101 = 10'h1d == addr; // @[Conditional.scala 37:30:@2147.62]
  assign _T_104 = 10'h1e == addr; // @[Conditional.scala 37:30:@2152.64]
  assign _T_107 = 10'h1f == addr; // @[Conditional.scala 37:30:@2157.66]
  assign _T_110 = 10'h20 == addr; // @[Conditional.scala 37:30:@2162.68]
  assign _T_113 = 10'h21 == addr; // @[Conditional.scala 37:30:@2167.70]
  assign _T_116 = 10'h22 == addr; // @[Conditional.scala 37:30:@2172.72]
  assign _T_119 = 10'h23 == addr; // @[Conditional.scala 37:30:@2177.74]
  assign _T_122 = 10'h24 == addr; // @[Conditional.scala 37:30:@2182.76]
  assign _T_125 = 10'h25 == addr; // @[Conditional.scala 37:30:@2187.78]
  assign _T_128 = 10'h26 == addr; // @[Conditional.scala 37:30:@2192.80]
  assign _T_131 = 10'h27 == addr; // @[Conditional.scala 37:30:@2197.82]
  assign _T_134 = 10'h28 == addr; // @[Conditional.scala 37:30:@2202.84]
  assign _T_137 = 10'h29 == addr; // @[Conditional.scala 37:30:@2207.86]
  assign _T_140 = 10'h2a == addr; // @[Conditional.scala 37:30:@2212.88]
  assign _T_143 = 10'h2b == addr; // @[Conditional.scala 37:30:@2217.90]
  assign _T_146 = 10'h2c == addr; // @[Conditional.scala 37:30:@2222.92]
  assign _T_149 = 10'h2d == addr; // @[Conditional.scala 37:30:@2227.94]
  assign _T_152 = 10'h2e == addr; // @[Conditional.scala 37:30:@2232.96]
  assign _T_155 = 10'h2f == addr; // @[Conditional.scala 37:30:@2237.98]
  assign _T_158 = 10'h30 == addr; // @[Conditional.scala 37:30:@2242.100]
  assign _T_161 = 10'h31 == addr; // @[Conditional.scala 37:30:@2247.102]
  assign _T_164 = 10'h32 == addr; // @[Conditional.scala 37:30:@2252.104]
  assign _T_167 = 10'h33 == addr; // @[Conditional.scala 37:30:@2257.106]
  assign _T_170 = 10'h34 == addr; // @[Conditional.scala 37:30:@2262.108]
  assign _T_173 = 10'h35 == addr; // @[Conditional.scala 37:30:@2267.110]
  assign _T_176 = 10'h36 == addr; // @[Conditional.scala 37:30:@2272.112]
  assign _T_179 = 10'h37 == addr; // @[Conditional.scala 37:30:@2277.114]
  assign _T_182 = 10'h38 == addr; // @[Conditional.scala 37:30:@2282.116]
  assign _T_185 = 10'h39 == addr; // @[Conditional.scala 37:30:@2287.118]
  assign _T_188 = 10'h3a == addr; // @[Conditional.scala 37:30:@2292.120]
  assign _T_191 = 10'h3b == addr; // @[Conditional.scala 37:30:@2297.122]
  assign _T_194 = 10'h3c == addr; // @[Conditional.scala 37:30:@2302.124]
  assign _T_197 = 10'h3d == addr; // @[Conditional.scala 37:30:@2307.126]
  assign _T_200 = 10'h3e == addr; // @[Conditional.scala 37:30:@2312.128]
  assign _T_203 = 10'h3f == addr; // @[Conditional.scala 37:30:@2317.130]
  assign _T_206 = 10'h40 == addr; // @[Conditional.scala 37:30:@2322.132]
  assign _T_209 = 10'h41 == addr; // @[Conditional.scala 37:30:@2327.134]
  assign _T_212 = 10'h42 == addr; // @[Conditional.scala 37:30:@2332.136]
  assign _T_215 = 10'h43 == addr; // @[Conditional.scala 37:30:@2337.138]
  assign _T_218 = 10'h44 == addr; // @[Conditional.scala 37:30:@2342.140]
  assign _T_221 = 10'h45 == addr; // @[Conditional.scala 37:30:@2347.142]
  assign _T_224 = 10'h46 == addr; // @[Conditional.scala 37:30:@2352.144]
  assign _T_227 = 10'h47 == addr; // @[Conditional.scala 37:30:@2357.146]
  assign _T_230 = 10'h48 == addr; // @[Conditional.scala 37:30:@2362.148]
  assign _T_233 = 10'h49 == addr; // @[Conditional.scala 37:30:@2367.150]
  assign _T_236 = 10'h4a == addr; // @[Conditional.scala 37:30:@2372.152]
  assign _T_239 = 10'h4b == addr; // @[Conditional.scala 37:30:@2377.154]
  assign _T_242 = 10'h4c == addr; // @[Conditional.scala 37:30:@2382.156]
  assign _T_245 = 10'h4d == addr; // @[Conditional.scala 37:30:@2387.158]
  assign _T_248 = 10'h4e == addr; // @[Conditional.scala 37:30:@2392.160]
  assign _T_251 = 10'h4f == addr; // @[Conditional.scala 37:30:@2397.162]
  assign _T_254 = 10'h50 == addr; // @[Conditional.scala 37:30:@2402.164]
  assign _T_257 = 10'h51 == addr; // @[Conditional.scala 37:30:@2407.166]
  assign _T_260 = 10'h52 == addr; // @[Conditional.scala 37:30:@2412.168]
  assign _T_263 = 10'h53 == addr; // @[Conditional.scala 37:30:@2417.170]
  assign _T_266 = 10'h54 == addr; // @[Conditional.scala 37:30:@2422.172]
  assign _T_269 = 10'h55 == addr; // @[Conditional.scala 37:30:@2427.174]
  assign _T_272 = 10'h56 == addr; // @[Conditional.scala 37:30:@2432.176]
  assign _T_275 = 10'h57 == addr; // @[Conditional.scala 37:30:@2437.178]
  assign _T_278 = 10'h58 == addr; // @[Conditional.scala 37:30:@2442.180]
  assign _T_281 = 10'h59 == addr; // @[Conditional.scala 37:30:@2447.182]
  assign _T_284 = 10'h5a == addr; // @[Conditional.scala 37:30:@2452.184]
  assign _T_287 = 10'h5b == addr; // @[Conditional.scala 37:30:@2457.186]
  assign _T_290 = 10'h5c == addr; // @[Conditional.scala 37:30:@2462.188]
  assign _T_293 = 10'h5d == addr; // @[Conditional.scala 37:30:@2467.190]
  assign _T_296 = 10'h5e == addr; // @[Conditional.scala 37:30:@2472.192]
  assign _T_299 = 10'h5f == addr; // @[Conditional.scala 37:30:@2477.194]
  assign _T_302 = 10'h60 == addr; // @[Conditional.scala 37:30:@2482.196]
  assign _T_305 = 10'h61 == addr; // @[Conditional.scala 37:30:@2487.198]
  assign _T_308 = 10'h62 == addr; // @[Conditional.scala 37:30:@2492.200]
  assign _T_311 = 10'h63 == addr; // @[Conditional.scala 37:30:@2497.202]
  assign _T_314 = 10'h64 == addr; // @[Conditional.scala 37:30:@2502.204]
  assign _T_317 = 10'h65 == addr; // @[Conditional.scala 37:30:@2507.206]
  assign _T_320 = 10'h66 == addr; // @[Conditional.scala 37:30:@2512.208]
  assign _T_323 = 10'h67 == addr; // @[Conditional.scala 37:30:@2517.210]
  assign _T_326 = 10'h68 == addr; // @[Conditional.scala 37:30:@2522.212]
  assign _T_329 = 10'h69 == addr; // @[Conditional.scala 37:30:@2527.214]
  assign _T_332 = 10'h6a == addr; // @[Conditional.scala 37:30:@2532.216]
  assign _T_335 = 10'h6b == addr; // @[Conditional.scala 37:30:@2537.218]
  assign _T_338 = 10'h6c == addr; // @[Conditional.scala 37:30:@2542.220]
  assign _T_341 = 10'h6d == addr; // @[Conditional.scala 37:30:@2547.222]
  assign _T_344 = 10'h6e == addr; // @[Conditional.scala 37:30:@2552.224]
  assign _T_347 = 10'h6f == addr; // @[Conditional.scala 37:30:@2557.226]
  assign _T_350 = 10'h70 == addr; // @[Conditional.scala 37:30:@2562.228]
  assign _T_353 = 10'h71 == addr; // @[Conditional.scala 37:30:@2567.230]
  assign _T_356 = 10'h72 == addr; // @[Conditional.scala 37:30:@2572.232]
  assign _T_359 = 10'h73 == addr; // @[Conditional.scala 37:30:@2577.234]
  assign _T_362 = 10'h74 == addr; // @[Conditional.scala 37:30:@2582.236]
  assign _T_365 = 10'h75 == addr; // @[Conditional.scala 37:30:@2587.238]
  assign _T_368 = 10'h76 == addr; // @[Conditional.scala 37:30:@2592.240]
  assign _T_371 = 10'h77 == addr; // @[Conditional.scala 37:30:@2597.242]
  assign _T_374 = 10'h78 == addr; // @[Conditional.scala 37:30:@2602.244]
  assign _T_377 = 10'h79 == addr; // @[Conditional.scala 37:30:@2607.246]
  assign _T_380 = 10'h7a == addr; // @[Conditional.scala 37:30:@2612.248]
  assign _T_383 = 10'h7b == addr; // @[Conditional.scala 37:30:@2617.250]
  assign _T_386 = 10'h7c == addr; // @[Conditional.scala 37:30:@2622.252]
  assign _T_389 = 10'h7d == addr; // @[Conditional.scala 37:30:@2627.254]
  assign _T_392 = 10'h7e == addr; // @[Conditional.scala 37:30:@2632.256]
  assign _T_395 = 10'h7f == addr; // @[Conditional.scala 37:30:@2637.258]
  assign _T_398 = 10'h80 == addr; // @[Conditional.scala 37:30:@2642.260]
  assign _T_401 = 10'h81 == addr; // @[Conditional.scala 37:30:@2647.262]
  assign _T_404 = 10'h82 == addr; // @[Conditional.scala 37:30:@2652.264]
  assign _T_407 = 10'h83 == addr; // @[Conditional.scala 37:30:@2657.266]
  assign _T_410 = 10'h84 == addr; // @[Conditional.scala 37:30:@2662.268]
  assign _T_413 = 10'h85 == addr; // @[Conditional.scala 37:30:@2667.270]
  assign _T_416 = 10'h86 == addr; // @[Conditional.scala 37:30:@2672.272]
  assign _T_419 = 10'h87 == addr; // @[Conditional.scala 37:30:@2677.274]
  assign _T_422 = 10'h88 == addr; // @[Conditional.scala 37:30:@2682.276]
  assign _T_425 = 10'h89 == addr; // @[Conditional.scala 37:30:@2687.278]
  assign _T_428 = 10'h8a == addr; // @[Conditional.scala 37:30:@2692.280]
  assign _T_431 = 10'h8b == addr; // @[Conditional.scala 37:30:@2697.282]
  assign _T_434 = 10'h8c == addr; // @[Conditional.scala 37:30:@2702.284]
  assign _T_437 = 10'h8d == addr; // @[Conditional.scala 37:30:@2707.286]
  assign _T_440 = 10'h8e == addr; // @[Conditional.scala 37:30:@2712.288]
  assign _T_443 = 10'h8f == addr; // @[Conditional.scala 37:30:@2717.290]
  assign _T_446 = 10'h90 == addr; // @[Conditional.scala 37:30:@2722.292]
  assign _T_449 = 10'h91 == addr; // @[Conditional.scala 37:30:@2727.294]
  assign _T_452 = 10'h92 == addr; // @[Conditional.scala 37:30:@2732.296]
  assign _T_455 = 10'h93 == addr; // @[Conditional.scala 37:30:@2737.298]
  assign _T_458 = 10'h94 == addr; // @[Conditional.scala 37:30:@2742.300]
  assign _T_461 = 10'h95 == addr; // @[Conditional.scala 37:30:@2747.302]
  assign _T_464 = 10'h96 == addr; // @[Conditional.scala 37:30:@2752.304]
  assign _T_467 = 10'h97 == addr; // @[Conditional.scala 37:30:@2757.306]
  assign _T_470 = 10'h98 == addr; // @[Conditional.scala 37:30:@2762.308]
  assign _T_473 = 10'h99 == addr; // @[Conditional.scala 37:30:@2767.310]
  assign _T_476 = 10'h9a == addr; // @[Conditional.scala 37:30:@2772.312]
  assign _T_479 = 10'h9b == addr; // @[Conditional.scala 37:30:@2777.314]
  assign _T_482 = 10'h9c == addr; // @[Conditional.scala 37:30:@2782.316]
  assign _T_485 = 10'h9d == addr; // @[Conditional.scala 37:30:@2787.318]
  assign _T_488 = 10'h9e == addr; // @[Conditional.scala 37:30:@2792.320]
  assign _T_491 = 10'h9f == addr; // @[Conditional.scala 37:30:@2797.322]
  assign _T_494 = 10'ha0 == addr; // @[Conditional.scala 37:30:@2802.324]
  assign _T_497 = 10'ha1 == addr; // @[Conditional.scala 37:30:@2807.326]
  assign _T_500 = 10'ha2 == addr; // @[Conditional.scala 37:30:@2812.328]
  assign _T_503 = 10'ha3 == addr; // @[Conditional.scala 37:30:@2817.330]
  assign _T_506 = 10'ha4 == addr; // @[Conditional.scala 37:30:@2822.332]
  assign _T_509 = 10'ha5 == addr; // @[Conditional.scala 37:30:@2827.334]
  assign _T_512 = 10'ha6 == addr; // @[Conditional.scala 37:30:@2832.336]
  assign _T_515 = 10'ha7 == addr; // @[Conditional.scala 37:30:@2837.338]
  assign _T_518 = 10'ha8 == addr; // @[Conditional.scala 37:30:@2842.340]
  assign _T_521 = 10'ha9 == addr; // @[Conditional.scala 37:30:@2847.342]
  assign _T_524 = 10'haa == addr; // @[Conditional.scala 37:30:@2852.344]
  assign _T_527 = 10'hab == addr; // @[Conditional.scala 37:30:@2857.346]
  assign _T_530 = 10'hac == addr; // @[Conditional.scala 37:30:@2862.348]
  assign _T_533 = 10'had == addr; // @[Conditional.scala 37:30:@2867.350]
  assign _T_536 = 10'hae == addr; // @[Conditional.scala 37:30:@2872.352]
  assign _T_539 = 10'haf == addr; // @[Conditional.scala 37:30:@2877.354]
  assign _T_542 = 10'hb0 == addr; // @[Conditional.scala 37:30:@2882.356]
  assign _T_545 = 10'hb1 == addr; // @[Conditional.scala 37:30:@2887.358]
  assign _T_548 = 10'hb2 == addr; // @[Conditional.scala 37:30:@2892.360]
  assign _T_551 = 10'hb3 == addr; // @[Conditional.scala 37:30:@2897.362]
  assign _T_554 = 10'hb4 == addr; // @[Conditional.scala 37:30:@2902.364]
  assign _T_557 = 10'hb5 == addr; // @[Conditional.scala 37:30:@2907.366]
  assign _T_560 = 10'hb6 == addr; // @[Conditional.scala 37:30:@2912.368]
  assign _T_563 = 10'hb7 == addr; // @[Conditional.scala 37:30:@2917.370]
  assign _T_566 = 10'hb8 == addr; // @[Conditional.scala 37:30:@2922.372]
  assign _T_569 = 10'hb9 == addr; // @[Conditional.scala 37:30:@2927.374]
  assign _T_572 = 10'hba == addr; // @[Conditional.scala 37:30:@2932.376]
  assign _T_575 = 10'hbb == addr; // @[Conditional.scala 37:30:@2937.378]
  assign _T_578 = 10'hbc == addr; // @[Conditional.scala 37:30:@2942.380]
  assign _T_581 = 10'hbd == addr; // @[Conditional.scala 37:30:@2947.382]
  assign _T_584 = 10'hbe == addr; // @[Conditional.scala 37:30:@2952.384]
  assign _T_587 = 10'hbf == addr; // @[Conditional.scala 37:30:@2957.386]
  assign _T_590 = 10'hc0 == addr; // @[Conditional.scala 37:30:@2962.388]
  assign _T_593 = 10'hc1 == addr; // @[Conditional.scala 37:30:@2967.390]
  assign _T_596 = 10'hc2 == addr; // @[Conditional.scala 37:30:@2972.392]
  assign _T_599 = 10'hc3 == addr; // @[Conditional.scala 37:30:@2977.394]
  assign _T_602 = 10'hc4 == addr; // @[Conditional.scala 37:30:@2982.396]
  assign _T_605 = 10'hc5 == addr; // @[Conditional.scala 37:30:@2987.398]
  assign _T_608 = 10'hc6 == addr; // @[Conditional.scala 37:30:@2992.400]
  assign _T_611 = 10'hc7 == addr; // @[Conditional.scala 37:30:@2997.402]
  assign _T_614 = 10'hc8 == addr; // @[Conditional.scala 37:30:@3002.404]
  assign _T_617 = 10'hc9 == addr; // @[Conditional.scala 37:30:@3007.406]
  assign _T_620 = 10'hca == addr; // @[Conditional.scala 37:30:@3012.408]
  assign _T_623 = 10'hcb == addr; // @[Conditional.scala 37:30:@3017.410]
  assign _T_626 = 10'hcc == addr; // @[Conditional.scala 37:30:@3022.412]
  assign _T_629 = 10'hcd == addr; // @[Conditional.scala 37:30:@3027.414]
  assign _T_632 = 10'hce == addr; // @[Conditional.scala 37:30:@3032.416]
  assign _T_635 = 10'hcf == addr; // @[Conditional.scala 37:30:@3037.418]
  assign _T_638 = 10'hd0 == addr; // @[Conditional.scala 37:30:@3042.420]
  assign _T_641 = 10'hd1 == addr; // @[Conditional.scala 37:30:@3047.422]
  assign _T_644 = 10'hd2 == addr; // @[Conditional.scala 37:30:@3052.424]
  assign _T_647 = 10'hd3 == addr; // @[Conditional.scala 37:30:@3057.426]
  assign _T_650 = 10'hd4 == addr; // @[Conditional.scala 37:30:@3062.428]
  assign _T_653 = 10'hd5 == addr; // @[Conditional.scala 37:30:@3067.430]
  assign _T_656 = 10'hd6 == addr; // @[Conditional.scala 37:30:@3072.432]
  assign _T_659 = 10'hd7 == addr; // @[Conditional.scala 37:30:@3077.434]
  assign _T_662 = 10'hd8 == addr; // @[Conditional.scala 37:30:@3082.436]
  assign _T_665 = 10'hd9 == addr; // @[Conditional.scala 37:30:@3087.438]
  assign _GEN_0 = _T_665 ? 32'h8067 : bmem_data; // @[Conditional.scala 39:67:@3088.438]
  assign _GEN_1 = _T_662 ? 32'h3010113 : _GEN_0; // @[Conditional.scala 39:67:@3083.436]
  assign _GEN_2 = _T_659 ? 32'h2812403 : _GEN_1; // @[Conditional.scala 39:67:@3078.434]
  assign _GEN_3 = _T_656 ? 32'h2c12083 : _GEN_2; // @[Conditional.scala 39:67:@3073.432]
  assign _GEN_4 = _T_653 ? 32'h13 : _GEN_3; // @[Conditional.scala 39:67:@3068.430]
  assign _GEN_5 = _T_650 ? 32'hfc07dce3 : _GEN_4; // @[Conditional.scala 39:67:@3063.428]
  assign _GEN_6 = _T_647 ? 32'hfec42783 : _GEN_5; // @[Conditional.scala 39:67:@3058.426]
  assign _GEN_7 = _T_644 ? 32'hfef42623 : _GEN_6; // @[Conditional.scala 39:67:@3053.424]
  assign _GEN_8 = _T_641 ? 32'hfff78793 : _GEN_7; // @[Conditional.scala 39:67:@3048.422]
  assign _GEN_9 = _T_638 ? 32'hfec42783 : _GEN_8; // @[Conditional.scala 39:67:@3043.420]
  assign _GEN_10 = _T_635 ? 32'hd25ff0ef : _GEN_9; // @[Conditional.scala 39:67:@3038.418]
  assign _GEN_11 = _T_632 ? 32'h78513 : _GEN_10; // @[Conditional.scala 39:67:@3033.416]
  assign _GEN_12 = _T_629 ? 32'hff87c783 : _GEN_11; // @[Conditional.scala 39:67:@3028.414]
  assign _GEN_13 = _T_626 ? 32'hf707b3 : _GEN_12; // @[Conditional.scala 39:67:@3023.412]
  assign _GEN_14 = _T_623 ? 32'hff040713 : _GEN_13; // @[Conditional.scala 39:67:@3018.410]
  assign _GEN_15 = _T_620 ? 32'hfec42783 : _GEN_14; // @[Conditional.scala 39:67:@3013.408]
  assign _GEN_16 = _T_617 ? 32'h280006f : _GEN_15; // @[Conditional.scala 39:67:@3008.406]
  assign _GEN_17 = _T_614 ? 32'hfef42623 : _GEN_16; // @[Conditional.scala 39:67:@3003.404]
  assign _GEN_18 = _T_611 ? 32'h200793 : _GEN_17; // @[Conditional.scala 39:67:@2998.402]
  assign _GEN_19 = _T_608 ? 32'hfef42423 : _GEN_18; // @[Conditional.scala 39:67:@2993.400]
  assign _GEN_20 = _T_605 ? 32'hfdc42783 : _GEN_19; // @[Conditional.scala 39:67:@2988.398]
  assign _GEN_21 = _T_602 ? 32'hfca42e23 : _GEN_20; // @[Conditional.scala 39:67:@2983.396]
  assign _GEN_22 = _T_599 ? 32'h3010413 : _GEN_21; // @[Conditional.scala 39:67:@2978.394]
  assign _GEN_23 = _T_596 ? 32'h2812423 : _GEN_22; // @[Conditional.scala 39:67:@2973.392]
  assign _GEN_24 = _T_593 ? 32'h2112623 : _GEN_23; // @[Conditional.scala 39:67:@2968.390]
  assign _GEN_25 = _T_590 ? 32'hfd010113 : _GEN_24; // @[Conditional.scala 39:67:@2963.388]
  assign _GEN_26 = _T_587 ? 32'h8067 : _GEN_25; // @[Conditional.scala 39:67:@2958.386]
  assign _GEN_27 = _T_584 ? 32'h3010113 : _GEN_26; // @[Conditional.scala 39:67:@2953.384]
  assign _GEN_28 = _T_581 ? 32'h2812403 : _GEN_27; // @[Conditional.scala 39:67:@2948.382]
  assign _GEN_29 = _T_578 ? 32'h2c12083 : _GEN_28; // @[Conditional.scala 39:67:@2943.380]
  assign _GEN_30 = _T_575 ? 32'h78513 : _GEN_29; // @[Conditional.scala 39:67:@2938.378]
  assign _GEN_31 = _T_572 ? 32'hfe842783 : _GEN_30; // @[Conditional.scala 39:67:@2933.376]
  assign _GEN_32 = _T_569 ? 32'he782a3 : _GEN_31; // @[Conditional.scala 39:67:@2928.374]
  assign _GEN_33 = _T_566 ? 32'hff77713 : _GEN_32; // @[Conditional.scala 39:67:@2923.372]
  assign _GEN_34 = _T_563 ? 32'hffe77713 : _GEN_33; // @[Conditional.scala 39:67:@2918.370]
  assign _GEN_35 = _T_560 ? 32'h37b7 : _GEN_34; // @[Conditional.scala 39:67:@2913.368]
  assign _GEN_36 = _T_557 ? 32'hff7f713 : _GEN_35; // @[Conditional.scala 39:67:@2908.366]
  assign _GEN_37 = _T_554 ? 32'h57c783 : _GEN_36; // @[Conditional.scala 39:67:@2903.364]
  assign _GEN_38 = _T_551 ? 32'h37b7 : _GEN_37; // @[Conditional.scala 39:67:@2898.362]
  assign _GEN_39 = _T_548 ? 32'hfce7f6e3 : _GEN_38; // @[Conditional.scala 39:67:@2893.360]
  assign _GEN_40 = _T_545 ? 32'h300793 : _GEN_39; // @[Conditional.scala 39:67:@2888.358]
  assign _GEN_41 = _T_542 ? 32'hfec42703 : _GEN_40; // @[Conditional.scala 39:67:@2883.356]
  assign _GEN_42 = _T_539 ? 32'hfef42623 : _GEN_41; // @[Conditional.scala 39:67:@2878.354]
  assign _GEN_43 = _T_536 ? 32'h178793 : _GEN_42; // @[Conditional.scala 39:67:@2873.352]
  assign _GEN_44 = _T_533 ? 32'hfec42783 : _GEN_43; // @[Conditional.scala 39:67:@2868.350]
  assign _GEN_45 = _T_530 ? 32'hfee78c23 : _GEN_44; // @[Conditional.scala 39:67:@2863.348]
  assign _GEN_46 = _T_527 ? 32'hf687b3 : _GEN_45; // @[Conditional.scala 39:67:@2858.346]
  assign _GEN_47 = _T_524 ? 32'hff040693 : _GEN_46; // @[Conditional.scala 39:67:@2853.344]
  assign _GEN_48 = _T_521 ? 32'hfec42783 : _GEN_47; // @[Conditional.scala 39:67:@2848.342]
  assign _GEN_49 = _T_518 ? 32'h78713 : _GEN_48; // @[Conditional.scala 39:67:@2843.340]
  assign _GEN_50 = _T_515 ? 32'h50793 : _GEN_49; // @[Conditional.scala 39:67:@2838.338]
  assign _GEN_51 = _T_512 ? 32'hdc9ff0ef : _GEN_50; // @[Conditional.scala 39:67:@2833.336]
  assign _GEN_52 = _T_509 ? 32'h513 : _GEN_51; // @[Conditional.scala 39:67:@2828.334]
  assign _GEN_53 = _T_506 ? 32'h300006f : _GEN_52; // @[Conditional.scala 39:67:@2823.332]
  assign _GEN_54 = _T_503 ? 32'hfe042623 : _GEN_53; // @[Conditional.scala 39:67:@2818.330]
  assign _GEN_55 = _T_500 ? 32'h78000ef : _GEN_54; // @[Conditional.scala 39:67:@2813.328]
  assign _GEN_56 = _T_497 ? 32'hfdc42503 : _GEN_55; // @[Conditional.scala 39:67:@2808.326]
  assign _GEN_57 = _T_494 ? 32'hde1ff0ef : _GEN_56; // @[Conditional.scala 39:67:@2803.324]
  assign _GEN_58 = _T_491 ? 32'h300513 : _GEN_57; // @[Conditional.scala 39:67:@2798.322]
  assign _GEN_59 = _T_488 ? 32'he782a3 : _GEN_58; // @[Conditional.scala 39:67:@2793.320]
  assign _GEN_60 = _T_485 ? 32'hff77713 : _GEN_59; // @[Conditional.scala 39:67:@2788.318]
  assign _GEN_61 = _T_482 ? 32'h176713 : _GEN_60; // @[Conditional.scala 39:67:@2783.316]
  assign _GEN_62 = _T_479 ? 32'h37b7 : _GEN_61; // @[Conditional.scala 39:67:@2778.314]
  assign _GEN_63 = _T_476 ? 32'hff7f713 : _GEN_62; // @[Conditional.scala 39:67:@2773.312]
  assign _GEN_64 = _T_473 ? 32'h57c783 : _GEN_63; // @[Conditional.scala 39:67:@2768.310]
  assign _GEN_65 = _T_470 ? 32'h37b7 : _GEN_64; // @[Conditional.scala 39:67:@2763.308]
  assign _GEN_66 = _T_467 ? 32'hfca42e23 : _GEN_65; // @[Conditional.scala 39:67:@2758.306]
  assign _GEN_67 = _T_464 ? 32'h3010413 : _GEN_66; // @[Conditional.scala 39:67:@2753.304]
  assign _GEN_68 = _T_461 ? 32'h2812423 : _GEN_67; // @[Conditional.scala 39:67:@2748.302]
  assign _GEN_69 = _T_458 ? 32'h2112623 : _GEN_68; // @[Conditional.scala 39:67:@2743.300]
  assign _GEN_70 = _T_455 ? 32'hfd010113 : _GEN_69; // @[Conditional.scala 39:67:@2738.298]
  assign _GEN_71 = _T_452 ? 32'h8067 : _GEN_70; // @[Conditional.scala 39:67:@2733.296]
  assign _GEN_72 = _T_449 ? 32'h3010113 : _GEN_71; // @[Conditional.scala 39:67:@2728.294]
  assign _GEN_73 = _T_446 ? 32'h2812403 : _GEN_72; // @[Conditional.scala 39:67:@2723.292]
  assign _GEN_74 = _T_443 ? 32'h2c12083 : _GEN_73; // @[Conditional.scala 39:67:@2718.290]
  assign _GEN_75 = _T_440 ? 32'h13 : _GEN_74; // @[Conditional.scala 39:67:@2713.288]
  assign _GEN_76 = _T_437 ? 32'hfaf76ee3 : _GEN_75; // @[Conditional.scala 39:67:@2708.286]
  assign _GEN_77 = _T_434 ? 32'hfe842703 : _GEN_76; // @[Conditional.scala 39:67:@2703.284]
  assign _GEN_78 = _T_431 ? 32'h27d793 : _GEN_77; // @[Conditional.scala 39:67:@2698.282]
  assign _GEN_79 = _T_428 ? 32'hfe042783 : _GEN_78; // @[Conditional.scala 39:67:@2693.280]
  assign _GEN_80 = _T_425 ? 32'hfef42623 : _GEN_79; // @[Conditional.scala 39:67:@2688.278]
  assign _GEN_81 = _T_422 ? 32'h478793 : _GEN_80; // @[Conditional.scala 39:67:@2683.276]
  assign _GEN_82 = _T_419 ? 32'hfec42783 : _GEN_81; // @[Conditional.scala 39:67:@2678.274]
  assign _GEN_83 = _T_416 ? 32'he7a023 : _GEN_82; // @[Conditional.scala 39:67:@2673.272]
  assign _GEN_84 = _T_413 ? 32'hfd842703 : _GEN_83; // @[Conditional.scala 39:67:@2668.270]
  assign _GEN_85 = _T_410 ? 32'hf707b3 : _GEN_84; // @[Conditional.scala 39:67:@2663.268]
  assign _GEN_86 = _T_407 ? 32'hfdc42703 : _GEN_85; // @[Conditional.scala 39:67:@2658.266]
  assign _GEN_87 = _T_404 ? 32'h279793 : _GEN_86; // @[Conditional.scala 39:67:@2653.264]
  assign _GEN_88 = _T_401 ? 32'hfee42423 : _GEN_87; // @[Conditional.scala 39:67:@2648.262]
  assign _GEN_89 = _T_398 ? 32'h178713 : _GEN_88; // @[Conditional.scala 39:67:@2643.260]
  assign _GEN_90 = _T_395 ? 32'hfe842783 : _GEN_89; // @[Conditional.scala 39:67:@2638.258]
  assign _GEN_91 = _T_392 ? 32'hfca42c23 : _GEN_90; // @[Conditional.scala 39:67:@2633.256]
  assign _GEN_92 = _T_389 ? 32'h58000ef : _GEN_91; // @[Conditional.scala 39:67:@2628.254]
  assign _GEN_93 = _T_386 ? 32'hfec42503 : _GEN_92; // @[Conditional.scala 39:67:@2623.252]
  assign _GEN_94 = _T_383 ? 32'h3c0006f : _GEN_93; // @[Conditional.scala 39:67:@2618.250]
  assign _GEN_95 = _T_380 ? 32'hfef42623 : _GEN_94; // @[Conditional.scala 39:67:@2613.248]
  assign _GEN_96 = _T_377 ? 32'hc78793 : _GEN_95; // @[Conditional.scala 39:67:@2608.246]
  assign _GEN_97 = _T_374 ? 32'hfec42783 : _GEN_96; // @[Conditional.scala 39:67:@2603.244]
  assign _GEN_98 = _T_371 ? 32'hfe042423 : _GEN_97; // @[Conditional.scala 39:67:@2598.242]
  assign _GEN_99 = _T_368 ? 32'hfc042c23 : _GEN_98; // @[Conditional.scala 39:67:@2593.240]
  assign _GEN_100 = _T_365 ? 32'hfc042e23 : _GEN_99; // @[Conditional.scala 39:67:@2588.238]
  assign _GEN_101 = _T_362 ? 32'hfea42023 : _GEN_100; // @[Conditional.scala 39:67:@2583.236]
  assign _GEN_102 = _T_359 ? 32'h80000ef : _GEN_101; // @[Conditional.scala 39:67:@2578.234]
  assign _GEN_103 = _T_356 ? 32'h78513 : _GEN_102; // @[Conditional.scala 39:67:@2573.232]
  assign _GEN_104 = _T_353 ? 32'h478793 : _GEN_103; // @[Conditional.scala 39:67:@2568.230]
  assign _GEN_105 = _T_350 ? 32'hfec42783 : _GEN_104; // @[Conditional.scala 39:67:@2563.228]
  assign _GEN_106 = _T_347 ? 32'hfea42223 : _GEN_105; // @[Conditional.scala 39:67:@2558.226]
  assign _GEN_107 = _T_344 ? 32'h94000ef : _GEN_106; // @[Conditional.scala 39:67:@2553.224]
  assign _GEN_108 = _T_341 ? 32'hfec42503 : _GEN_107; // @[Conditional.scala 39:67:@2548.222]
  assign _GEN_109 = _T_338 ? 32'hfe042623 : _GEN_108; // @[Conditional.scala 39:67:@2543.220]
  assign _GEN_110 = _T_335 ? 32'h3010413 : _GEN_109; // @[Conditional.scala 39:67:@2538.218]
  assign _GEN_111 = _T_332 ? 32'h2812423 : _GEN_110; // @[Conditional.scala 39:67:@2533.216]
  assign _GEN_112 = _T_329 ? 32'h2112623 : _GEN_111; // @[Conditional.scala 39:67:@2528.214]
  assign _GEN_113 = _T_326 ? 32'hfd010113 : _GEN_112; // @[Conditional.scala 39:67:@2523.212]
  assign _GEN_114 = _T_323 ? 32'h8067 : _GEN_113; // @[Conditional.scala 39:67:@2518.210]
  assign _GEN_115 = _T_320 ? 32'h1010113 : _GEN_114; // @[Conditional.scala 39:67:@2513.208]
  assign _GEN_116 = _T_317 ? 32'hc12403 : _GEN_115; // @[Conditional.scala 39:67:@2508.206]
  assign _GEN_117 = _T_314 ? 32'h13 : _GEN_116; // @[Conditional.scala 39:67:@2503.204]
  assign _GEN_118 = _T_311 ? 32'h28067 : _GEN_117; // @[Conditional.scala 39:67:@2498.202]
  assign _GEN_119 = _T_308 ? 32'h2b7 : _GEN_118; // @[Conditional.scala 39:67:@2493.200]
  assign _GEN_120 = _T_305 ? 32'h1010413 : _GEN_119; // @[Conditional.scala 39:67:@2488.198]
  assign _GEN_121 = _T_302 ? 32'h812623 : _GEN_120; // @[Conditional.scala 39:67:@2483.196]
  assign _GEN_122 = _T_299 ? 32'hff010113 : _GEN_121; // @[Conditional.scala 39:67:@2478.194]
  assign _GEN_123 = _T_296 ? 32'h8067 : _GEN_122; // @[Conditional.scala 39:67:@2473.192]
  assign _GEN_124 = _T_293 ? 32'h1010113 : _GEN_123; // @[Conditional.scala 39:67:@2468.190]
  assign _GEN_125 = _T_290 ? 32'h812403 : _GEN_124; // @[Conditional.scala 39:67:@2463.188]
  assign _GEN_126 = _T_287 ? 32'hc12083 : _GEN_125; // @[Conditional.scala 39:67:@2458.186]
  assign _GEN_127 = _T_284 ? 32'h78513 : _GEN_126; // @[Conditional.scala 39:67:@2453.184]
  assign _GEN_128 = _T_281 ? 32'h793 : _GEN_127; // @[Conditional.scala 39:67:@2448.182]
  assign _GEN_129 = _T_278 ? 32'h1c000ef : _GEN_128; // @[Conditional.scala 39:67:@2443.180]
  assign _GEN_130 = _T_275 ? 32'hf89ff0ef : _GEN_129; // @[Conditional.scala 39:67:@2438.178]
  assign _GEN_131 = _T_272 ? 32'h6b00513 : _GEN_130; // @[Conditional.scala 39:67:@2433.176]
  assign _GEN_132 = _T_269 ? 32'hf91ff0ef : _GEN_131; // @[Conditional.scala 39:67:@2428.174]
  assign _GEN_133 = _T_266 ? 32'h4f00513 : _GEN_132; // @[Conditional.scala 39:67:@2423.172]
  assign _GEN_134 = _T_263 ? 32'h54000ef : _GEN_133; // @[Conditional.scala 39:67:@2418.170]
  assign _GEN_135 = _T_260 ? 32'hed5ff0ef : _GEN_134; // @[Conditional.scala 39:67:@2413.168]
  assign _GEN_136 = _T_257 ? 32'h800513 : _GEN_135; // @[Conditional.scala 39:67:@2408.166]
  assign _GEN_137 = _T_254 ? 32'hf75ff0ef : _GEN_136; // @[Conditional.scala 39:67:@2403.164]
  assign _GEN_138 = _T_251 ? 32'h1000513 : _GEN_137; // @[Conditional.scala 39:67:@2398.162]
  assign _GEN_139 = _T_248 ? 32'h1010413 : _GEN_138; // @[Conditional.scala 39:67:@2393.160]
  assign _GEN_140 = _T_245 ? 32'h812423 : _GEN_139; // @[Conditional.scala 39:67:@2388.158]
  assign _GEN_141 = _T_242 ? 32'h112623 : _GEN_140; // @[Conditional.scala 39:67:@2383.156]
  assign _GEN_142 = _T_239 ? 32'hff010113 : _GEN_141; // @[Conditional.scala 39:67:@2378.154]
  assign _GEN_143 = _T_236 ? 32'h8067 : _GEN_142; // @[Conditional.scala 39:67:@2373.152]
  assign _GEN_144 = _T_233 ? 32'h2010113 : _GEN_143; // @[Conditional.scala 39:67:@2368.150]
  assign _GEN_145 = _T_230 ? 32'h1c12403 : _GEN_144; // @[Conditional.scala 39:67:@2363.148]
  assign _GEN_146 = _T_227 ? 32'h13 : _GEN_145; // @[Conditional.scala 39:67:@2358.146]
  assign _GEN_147 = _T_224 ? 32'he780a3 : _GEN_146; // @[Conditional.scala 39:67:@2353.144]
  assign _GEN_148 = _T_221 ? 32'hfef44703 : _GEN_147; // @[Conditional.scala 39:67:@2348.142]
  assign _GEN_149 = _T_218 ? 32'h27b7 : _GEN_148; // @[Conditional.scala 39:67:@2343.140]
  assign _GEN_150 = _T_215 ? 32'hfe0788e3 : _GEN_149; // @[Conditional.scala 39:67:@2338.138]
  assign _GEN_151 = _T_212 ? 32'h27f793 : _GEN_150; // @[Conditional.scala 39:67:@2333.136]
  assign _GEN_152 = _T_209 ? 32'hff7f793 : _GEN_151; // @[Conditional.scala 39:67:@2328.134]
  assign _GEN_153 = _T_206 ? 32'h47c783 : _GEN_152; // @[Conditional.scala 39:67:@2323.132]
  assign _GEN_154 = _T_203 ? 32'h27b7 : _GEN_153; // @[Conditional.scala 39:67:@2318.130]
  assign _GEN_155 = _T_200 ? 32'h13 : _GEN_154; // @[Conditional.scala 39:67:@2313.128]
  assign _GEN_156 = _T_197 ? 32'hfef407a3 : _GEN_155; // @[Conditional.scala 39:67:@2308.126]
  assign _GEN_157 = _T_194 ? 32'h50793 : _GEN_156; // @[Conditional.scala 39:67:@2303.124]
  assign _GEN_158 = _T_191 ? 32'h2010413 : _GEN_157; // @[Conditional.scala 39:67:@2298.122]
  assign _GEN_159 = _T_188 ? 32'h812e23 : _GEN_158; // @[Conditional.scala 39:67:@2293.120]
  assign _GEN_160 = _T_185 ? 32'hfe010113 : _GEN_159; // @[Conditional.scala 39:67:@2288.118]
  assign _GEN_161 = _T_182 ? 32'h8067 : _GEN_160; // @[Conditional.scala 39:67:@2283.116]
  assign _GEN_162 = _T_179 ? 32'h2010113 : _GEN_161; // @[Conditional.scala 39:67:@2278.114]
  assign _GEN_163 = _T_176 ? 32'h1c12403 : _GEN_162; // @[Conditional.scala 39:67:@2273.112]
  assign _GEN_164 = _T_173 ? 32'h13 : _GEN_163; // @[Conditional.scala 39:67:@2268.110]
  assign _GEN_165 = _T_170 ? 32'he78123 : _GEN_164; // @[Conditional.scala 39:67:@2263.108]
  assign _GEN_166 = _T_167 ? 32'hfef44703 : _GEN_165; // @[Conditional.scala 39:67:@2258.106]
  assign _GEN_167 = _T_164 ? 32'h27b7 : _GEN_166; // @[Conditional.scala 39:67:@2253.104]
  assign _GEN_168 = _T_161 ? 32'hfef407a3 : _GEN_167; // @[Conditional.scala 39:67:@2248.102]
  assign _GEN_169 = _T_158 ? 32'h50793 : _GEN_168; // @[Conditional.scala 39:67:@2243.100]
  assign _GEN_170 = _T_155 ? 32'h2010413 : _GEN_169; // @[Conditional.scala 39:67:@2238.98]
  assign _GEN_171 = _T_152 ? 32'h812e23 : _GEN_170; // @[Conditional.scala 39:67:@2233.96]
  assign _GEN_172 = _T_149 ? 32'hfe010113 : _GEN_171; // @[Conditional.scala 39:67:@2228.94]
  assign _GEN_173 = _T_146 ? 32'h8067 : _GEN_172; // @[Conditional.scala 39:67:@2223.92]
  assign _GEN_174 = _T_143 ? 32'h2010113 : _GEN_173; // @[Conditional.scala 39:67:@2218.90]
  assign _GEN_175 = _T_140 ? 32'h1c12403 : _GEN_174; // @[Conditional.scala 39:67:@2213.88]
  assign _GEN_176 = _T_137 ? 32'h78513 : _GEN_175; // @[Conditional.scala 39:67:@2208.86]
  assign _GEN_177 = _T_134 ? 32'hff7f793 : _GEN_176; // @[Conditional.scala 39:67:@2203.84]
  assign _GEN_178 = _T_131 ? 32'h7c783 : _GEN_177; // @[Conditional.scala 39:67:@2198.82]
  assign _GEN_179 = _T_128 ? 32'h37b7 : _GEN_178; // @[Conditional.scala 39:67:@2193.80]
  assign _GEN_180 = _T_125 ? 32'hfe0788e3 : _GEN_179; // @[Conditional.scala 39:67:@2188.78]
  assign _GEN_181 = _T_122 ? 32'h107f793 : _GEN_180; // @[Conditional.scala 39:67:@2183.76]
  assign _GEN_182 = _T_119 ? 32'hff7f793 : _GEN_181; // @[Conditional.scala 39:67:@2178.74]
  assign _GEN_183 = _T_116 ? 32'h47c783 : _GEN_182; // @[Conditional.scala 39:67:@2173.72]
  assign _GEN_184 = _T_113 ? 32'h37b7 : _GEN_183; // @[Conditional.scala 39:67:@2168.70]
  assign _GEN_185 = _T_110 ? 32'h13 : _GEN_184; // @[Conditional.scala 39:67:@2163.68]
  assign _GEN_186 = _T_107 ? 32'he780a3 : _GEN_185; // @[Conditional.scala 39:67:@2158.66]
  assign _GEN_187 = _T_104 ? 32'hfef44703 : _GEN_186; // @[Conditional.scala 39:67:@2153.64]
  assign _GEN_188 = _T_101 ? 32'h37b7 : _GEN_187; // @[Conditional.scala 39:67:@2148.62]
  assign _GEN_189 = _T_98 ? 32'hfef407a3 : _GEN_188; // @[Conditional.scala 39:67:@2143.60]
  assign _GEN_190 = _T_95 ? 32'h50793 : _GEN_189; // @[Conditional.scala 39:67:@2138.58]
  assign _GEN_191 = _T_92 ? 32'h2010413 : _GEN_190; // @[Conditional.scala 39:67:@2133.56]
  assign _GEN_192 = _T_89 ? 32'h812e23 : _GEN_191; // @[Conditional.scala 39:67:@2128.54]
  assign _GEN_193 = _T_86 ? 32'hfe010113 : _GEN_192; // @[Conditional.scala 39:67:@2123.52]
  assign _GEN_194 = _T_83 ? 32'h8067 : _GEN_193; // @[Conditional.scala 39:67:@2118.50]
  assign _GEN_195 = _T_80 ? 32'h2010113 : _GEN_194; // @[Conditional.scala 39:67:@2113.48]
  assign _GEN_196 = _T_77 ? 32'h1c12403 : _GEN_195; // @[Conditional.scala 39:67:@2108.46]
  assign _GEN_197 = _T_74 ? 32'h13 : _GEN_196; // @[Conditional.scala 39:67:@2103.44]
  assign _GEN_198 = _T_71 ? 32'he78123 : _GEN_197; // @[Conditional.scala 39:67:@2098.42]
  assign _GEN_199 = _T_68 ? 32'hff77713 : _GEN_198; // @[Conditional.scala 39:67:@2093.40]
  assign _GEN_200 = _T_65 ? 32'he6e733 : _GEN_199; // @[Conditional.scala 39:67:@2088.38]
  assign _GEN_201 = _T_62 ? 32'hfef44703 : _GEN_200; // @[Conditional.scala 39:67:@2083.36]
  assign _GEN_202 = _T_59 ? 32'h37b7 : _GEN_201; // @[Conditional.scala 39:67:@2078.34]
  assign _GEN_203 = _T_56 ? 32'hff7f693 : _GEN_202; // @[Conditional.scala 39:67:@2073.32]
  assign _GEN_204 = _T_53 ? 32'h27c783 : _GEN_203; // @[Conditional.scala 39:67:@2068.30]
  assign _GEN_205 = _T_50 ? 32'h37b7 : _GEN_204; // @[Conditional.scala 39:67:@2063.28]
  assign _GEN_206 = _T_47 ? 32'hfef407a3 : _GEN_205; // @[Conditional.scala 39:67:@2058.26]
  assign _GEN_207 = _T_44 ? 32'h50793 : _GEN_206; // @[Conditional.scala 39:67:@2053.24]
  assign _GEN_208 = _T_41 ? 32'h2010413 : _GEN_207; // @[Conditional.scala 39:67:@2048.22]
  assign _GEN_209 = _T_38 ? 32'h812e23 : _GEN_208; // @[Conditional.scala 39:67:@2043.20]
  assign _GEN_210 = _T_35 ? 32'hfe010113 : _GEN_209; // @[Conditional.scala 39:67:@2038.18]
  assign _GEN_211 = _T_32 ? 32'h114000ef : _GEN_210; // @[Conditional.scala 39:67:@2033.16]
  assign _GEN_212 = _T_29 ? 32'h593 : _GEN_211; // @[Conditional.scala 39:67:@2028.14]
  assign _GEN_213 = _T_26 ? 32'h513 : _GEN_212; // @[Conditional.scala 39:67:@2023.12]
  assign _GEN_214 = _T_23 ? 32'hff810113 : _GEN_213; // @[Conditional.scala 39:67:@2018.10]
  assign _GEN_215 = _T_20 ? 32'hffffb117 : _GEN_214; // @[Conditional.scala 39:67:@2013.8]
  assign _GEN_216 = _T_17 ? 32'h40006f : _GEN_215; // @[Conditional.scala 39:67:@2008.6]
  assign _GEN_217 = _T_14 ? 32'h13 : _GEN_216; // @[Conditional.scala 40:58:@2003.4]
  assign io_bmem_rdata = bmem_data; // @[BMEM.scala 248:17:@3091.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bmem_data = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      bmem_data <= 32'h0;
    end else begin
      if (_T_14) begin
        bmem_data <= 32'h13;
      end else begin
        if (_T_17) begin
          bmem_data <= 32'h40006f;
        end else begin
          if (_T_20) begin
            bmem_data <= 32'hffffb117;
          end else begin
            if (_T_23) begin
              bmem_data <= 32'hff810113;
            end else begin
              if (_T_26) begin
                bmem_data <= 32'h513;
              end else begin
                if (_T_29) begin
                  bmem_data <= 32'h593;
                end else begin
                  if (_T_32) begin
                    bmem_data <= 32'h114000ef;
                  end else begin
                    if (_T_35) begin
                      bmem_data <= 32'hfe010113;
                    end else begin
                      if (_T_38) begin
                        bmem_data <= 32'h812e23;
                      end else begin
                        if (_T_41) begin
                          bmem_data <= 32'h2010413;
                        end else begin
                          if (_T_44) begin
                            bmem_data <= 32'h50793;
                          end else begin
                            if (_T_47) begin
                              bmem_data <= 32'hfef407a3;
                            end else begin
                              if (_T_50) begin
                                bmem_data <= 32'h37b7;
                              end else begin
                                if (_T_53) begin
                                  bmem_data <= 32'h27c783;
                                end else begin
                                  if (_T_56) begin
                                    bmem_data <= 32'hff7f693;
                                  end else begin
                                    if (_T_59) begin
                                      bmem_data <= 32'h37b7;
                                    end else begin
                                      if (_T_62) begin
                                        bmem_data <= 32'hfef44703;
                                      end else begin
                                        if (_T_65) begin
                                          bmem_data <= 32'he6e733;
                                        end else begin
                                          if (_T_68) begin
                                            bmem_data <= 32'hff77713;
                                          end else begin
                                            if (_T_71) begin
                                              bmem_data <= 32'he78123;
                                            end else begin
                                              if (_T_74) begin
                                                bmem_data <= 32'h13;
                                              end else begin
                                                if (_T_77) begin
                                                  bmem_data <= 32'h1c12403;
                                                end else begin
                                                  if (_T_80) begin
                                                    bmem_data <= 32'h2010113;
                                                  end else begin
                                                    if (_T_83) begin
                                                      bmem_data <= 32'h8067;
                                                    end else begin
                                                      if (_T_86) begin
                                                        bmem_data <= 32'hfe010113;
                                                      end else begin
                                                        if (_T_89) begin
                                                          bmem_data <= 32'h812e23;
                                                        end else begin
                                                          if (_T_92) begin
                                                            bmem_data <= 32'h2010413;
                                                          end else begin
                                                            if (_T_95) begin
                                                              bmem_data <= 32'h50793;
                                                            end else begin
                                                              if (_T_98) begin
                                                                bmem_data <= 32'hfef407a3;
                                                              end else begin
                                                                if (_T_101) begin
                                                                  bmem_data <= 32'h37b7;
                                                                end else begin
                                                                  if (_T_104) begin
                                                                    bmem_data <= 32'hfef44703;
                                                                  end else begin
                                                                    if (_T_107) begin
                                                                      bmem_data <= 32'he780a3;
                                                                    end else begin
                                                                      if (_T_110) begin
                                                                        bmem_data <= 32'h13;
                                                                      end else begin
                                                                        if (_T_113) begin
                                                                          bmem_data <= 32'h37b7;
                                                                        end else begin
                                                                          if (_T_116) begin
                                                                            bmem_data <= 32'h47c783;
                                                                          end else begin
                                                                            if (_T_119) begin
                                                                              bmem_data <= 32'hff7f793;
                                                                            end else begin
                                                                              if (_T_122) begin
                                                                                bmem_data <= 32'h107f793;
                                                                              end else begin
                                                                                if (_T_125) begin
                                                                                  bmem_data <= 32'hfe0788e3;
                                                                                end else begin
                                                                                  if (_T_128) begin
                                                                                    bmem_data <= 32'h37b7;
                                                                                  end else begin
                                                                                    if (_T_131) begin
                                                                                      bmem_data <= 32'h7c783;
                                                                                    end else begin
                                                                                      if (_T_134) begin
                                                                                        bmem_data <= 32'hff7f793;
                                                                                      end else begin
                                                                                        if (_T_137) begin
                                                                                          bmem_data <= 32'h78513;
                                                                                        end else begin
                                                                                          if (_T_140) begin
                                                                                            bmem_data <= 32'h1c12403;
                                                                                          end else begin
                                                                                            if (_T_143) begin
                                                                                              bmem_data <= 32'h2010113;
                                                                                            end else begin
                                                                                              if (_T_146) begin
                                                                                                bmem_data <= 32'h8067;
                                                                                              end else begin
                                                                                                if (_T_149) begin
                                                                                                  bmem_data <= 32'hfe010113;
                                                                                                end else begin
                                                                                                  if (_T_152) begin
                                                                                                    bmem_data <= 32'h812e23;
                                                                                                  end else begin
                                                                                                    if (_T_155) begin
                                                                                                      bmem_data <= 32'h2010413;
                                                                                                    end else begin
                                                                                                      if (_T_158) begin
                                                                                                        bmem_data <= 32'h50793;
                                                                                                      end else begin
                                                                                                        if (_T_161) begin
                                                                                                          bmem_data <= 32'hfef407a3;
                                                                                                        end else begin
                                                                                                          if (_T_164) begin
                                                                                                            bmem_data <= 32'h27b7;
                                                                                                          end else begin
                                                                                                            if (_T_167) begin
                                                                                                              bmem_data <= 32'hfef44703;
                                                                                                            end else begin
                                                                                                              if (_T_170) begin
                                                                                                                bmem_data <= 32'he78123;
                                                                                                              end else begin
                                                                                                                if (_T_173) begin
                                                                                                                  bmem_data <= 32'h13;
                                                                                                                end else begin
                                                                                                                  if (_T_176) begin
                                                                                                                    bmem_data <= 32'h1c12403;
                                                                                                                  end else begin
                                                                                                                    if (_T_179) begin
                                                                                                                      bmem_data <= 32'h2010113;
                                                                                                                    end else begin
                                                                                                                      if (_T_182) begin
                                                                                                                        bmem_data <= 32'h8067;
                                                                                                                      end else begin
                                                                                                                        if (_T_185) begin
                                                                                                                          bmem_data <= 32'hfe010113;
                                                                                                                        end else begin
                                                                                                                          if (_T_188) begin
                                                                                                                            bmem_data <= 32'h812e23;
                                                                                                                          end else begin
                                                                                                                            if (_T_191) begin
                                                                                                                              bmem_data <= 32'h2010413;
                                                                                                                            end else begin
                                                                                                                              if (_T_194) begin
                                                                                                                                bmem_data <= 32'h50793;
                                                                                                                              end else begin
                                                                                                                                if (_T_197) begin
                                                                                                                                  bmem_data <= 32'hfef407a3;
                                                                                                                                end else begin
                                                                                                                                  if (_T_200) begin
                                                                                                                                    bmem_data <= 32'h13;
                                                                                                                                  end else begin
                                                                                                                                    if (_T_203) begin
                                                                                                                                      bmem_data <= 32'h27b7;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_206) begin
                                                                                                                                        bmem_data <= 32'h47c783;
                                                                                                                                      end else begin
                                                                                                                                        if (_T_209) begin
                                                                                                                                          bmem_data <= 32'hff7f793;
                                                                                                                                        end else begin
                                                                                                                                          if (_T_212) begin
                                                                                                                                            bmem_data <= 32'h27f793;
                                                                                                                                          end else begin
                                                                                                                                            if (_T_215) begin
                                                                                                                                              bmem_data <= 32'hfe0788e3;
                                                                                                                                            end else begin
                                                                                                                                              if (_T_218) begin
                                                                                                                                                bmem_data <= 32'h27b7;
                                                                                                                                              end else begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  bmem_data <= 32'hfef44703;
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_224) begin
                                                                                                                                                    bmem_data <= 32'he780a3;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_227) begin
                                                                                                                                                      bmem_data <= 32'h13;
                                                                                                                                                    end else begin
                                                                                                                                                      if (_T_230) begin
                                                                                                                                                        bmem_data <= 32'h1c12403;
                                                                                                                                                      end else begin
                                                                                                                                                        if (_T_233) begin
                                                                                                                                                          bmem_data <= 32'h2010113;
                                                                                                                                                        end else begin
                                                                                                                                                          if (_T_236) begin
                                                                                                                                                            bmem_data <= 32'h8067;
                                                                                                                                                          end else begin
                                                                                                                                                            if (_T_239) begin
                                                                                                                                                              bmem_data <= 32'hff010113;
                                                                                                                                                            end else begin
                                                                                                                                                              if (_T_242) begin
                                                                                                                                                                bmem_data <= 32'h112623;
                                                                                                                                                              end else begin
                                                                                                                                                                if (_T_245) begin
                                                                                                                                                                  bmem_data <= 32'h812423;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (_T_248) begin
                                                                                                                                                                    bmem_data <= 32'h1010413;
                                                                                                                                                                  end else begin
                                                                                                                                                                    if (_T_251) begin
                                                                                                                                                                      bmem_data <= 32'h1000513;
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (_T_254) begin
                                                                                                                                                                        bmem_data <= 32'hf75ff0ef;
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (_T_257) begin
                                                                                                                                                                          bmem_data <= 32'h800513;
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (_T_260) begin
                                                                                                                                                                            bmem_data <= 32'hed5ff0ef;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (_T_263) begin
                                                                                                                                                                              bmem_data <= 32'h54000ef;
                                                                                                                                                                            end else begin
                                                                                                                                                                              if (_T_266) begin
                                                                                                                                                                                bmem_data <= 32'h4f00513;
                                                                                                                                                                              end else begin
                                                                                                                                                                                if (_T_269) begin
                                                                                                                                                                                  bmem_data <= 32'hf91ff0ef;
                                                                                                                                                                                end else begin
                                                                                                                                                                                  if (_T_272) begin
                                                                                                                                                                                    bmem_data <= 32'h6b00513;
                                                                                                                                                                                  end else begin
                                                                                                                                                                                    if (_T_275) begin
                                                                                                                                                                                      bmem_data <= 32'hf89ff0ef;
                                                                                                                                                                                    end else begin
                                                                                                                                                                                      if (_T_278) begin
                                                                                                                                                                                        bmem_data <= 32'h1c000ef;
                                                                                                                                                                                      end else begin
                                                                                                                                                                                        if (_T_281) begin
                                                                                                                                                                                          bmem_data <= 32'h793;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                          if (_T_284) begin
                                                                                                                                                                                            bmem_data <= 32'h78513;
                                                                                                                                                                                          end else begin
                                                                                                                                                                                            if (_T_287) begin
                                                                                                                                                                                              bmem_data <= 32'hc12083;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                              if (_T_290) begin
                                                                                                                                                                                                bmem_data <= 32'h812403;
                                                                                                                                                                                              end else begin
                                                                                                                                                                                                if (_T_293) begin
                                                                                                                                                                                                  bmem_data <= 32'h1010113;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                  if (_T_296) begin
                                                                                                                                                                                                    bmem_data <= 32'h8067;
                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                    if (_T_299) begin
                                                                                                                                                                                                      bmem_data <= 32'hff010113;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                      if (_T_302) begin
                                                                                                                                                                                                        bmem_data <= 32'h812623;
                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                        if (_T_305) begin
                                                                                                                                                                                                          bmem_data <= 32'h1010413;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                          if (_T_308) begin
                                                                                                                                                                                                            bmem_data <= 32'h2b7;
                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                            if (_T_311) begin
                                                                                                                                                                                                              bmem_data <= 32'h28067;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                              if (_T_314) begin
                                                                                                                                                                                                                bmem_data <= 32'h13;
                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                if (_T_317) begin
                                                                                                                                                                                                                  bmem_data <= 32'hc12403;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                  if (_T_320) begin
                                                                                                                                                                                                                    bmem_data <= 32'h1010113;
                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                    if (_T_323) begin
                                                                                                                                                                                                                      bmem_data <= 32'h8067;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                      if (_T_326) begin
                                                                                                                                                                                                                        bmem_data <= 32'hfd010113;
                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                        if (_T_329) begin
                                                                                                                                                                                                                          bmem_data <= 32'h2112623;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                          if (_T_332) begin
                                                                                                                                                                                                                            bmem_data <= 32'h2812423;
                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                            if (_T_335) begin
                                                                                                                                                                                                                              bmem_data <= 32'h3010413;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                              if (_T_338) begin
                                                                                                                                                                                                                                bmem_data <= 32'hfe042623;
                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                if (_T_341) begin
                                                                                                                                                                                                                                  bmem_data <= 32'hfec42503;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                  if (_T_344) begin
                                                                                                                                                                                                                                    bmem_data <= 32'h94000ef;
                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                    if (_T_347) begin
                                                                                                                                                                                                                                      bmem_data <= 32'hfea42223;
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                      if (_T_350) begin
                                                                                                                                                                                                                                        bmem_data <= 32'hfec42783;
                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                        if (_T_353) begin
                                                                                                                                                                                                                                          bmem_data <= 32'h478793;
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                          if (_T_356) begin
                                                                                                                                                                                                                                            bmem_data <= 32'h78513;
                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                            if (_T_359) begin
                                                                                                                                                                                                                                              bmem_data <= 32'h80000ef;
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                              if (_T_362) begin
                                                                                                                                                                                                                                                bmem_data <= 32'hfea42023;
                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                if (_T_365) begin
                                                                                                                                                                                                                                                  bmem_data <= 32'hfc042e23;
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                  if (_T_368) begin
                                                                                                                                                                                                                                                    bmem_data <= 32'hfc042c23;
                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                    if (_T_371) begin
                                                                                                                                                                                                                                                      bmem_data <= 32'hfe042423;
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                      if (_T_374) begin
                                                                                                                                                                                                                                                        bmem_data <= 32'hfec42783;
                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                        if (_T_377) begin
                                                                                                                                                                                                                                                          bmem_data <= 32'hc78793;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                          if (_T_380) begin
                                                                                                                                                                                                                                                            bmem_data <= 32'hfef42623;
                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                            if (_T_383) begin
                                                                                                                                                                                                                                                              bmem_data <= 32'h3c0006f;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                              if (_T_386) begin
                                                                                                                                                                                                                                                                bmem_data <= 32'hfec42503;
                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                if (_T_389) begin
                                                                                                                                                                                                                                                                  bmem_data <= 32'h58000ef;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                  if (_T_392) begin
                                                                                                                                                                                                                                                                    bmem_data <= 32'hfca42c23;
                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                    if (_T_395) begin
                                                                                                                                                                                                                                                                      bmem_data <= 32'hfe842783;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                      if (_T_398) begin
                                                                                                                                                                                                                                                                        bmem_data <= 32'h178713;
                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                        if (_T_401) begin
                                                                                                                                                                                                                                                                          bmem_data <= 32'hfee42423;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                          if (_T_404) begin
                                                                                                                                                                                                                                                                            bmem_data <= 32'h279793;
                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                            if (_T_407) begin
                                                                                                                                                                                                                                                                              bmem_data <= 32'hfdc42703;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                              if (_T_410) begin
                                                                                                                                                                                                                                                                                bmem_data <= 32'hf707b3;
                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                if (_T_413) begin
                                                                                                                                                                                                                                                                                  bmem_data <= 32'hfd842703;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                  if (_T_416) begin
                                                                                                                                                                                                                                                                                    bmem_data <= 32'he7a023;
                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                    if (_T_419) begin
                                                                                                                                                                                                                                                                                      bmem_data <= 32'hfec42783;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                      if (_T_422) begin
                                                                                                                                                                                                                                                                                        bmem_data <= 32'h478793;
                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                        if (_T_425) begin
                                                                                                                                                                                                                                                                                          bmem_data <= 32'hfef42623;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                          if (_T_428) begin
                                                                                                                                                                                                                                                                                            bmem_data <= 32'hfe042783;
                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                            if (_T_431) begin
                                                                                                                                                                                                                                                                                              bmem_data <= 32'h27d793;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                              if (_T_434) begin
                                                                                                                                                                                                                                                                                                bmem_data <= 32'hfe842703;
                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                if (_T_437) begin
                                                                                                                                                                                                                                                                                                  bmem_data <= 32'hfaf76ee3;
                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                  if (_T_440) begin
                                                                                                                                                                                                                                                                                                    bmem_data <= 32'h13;
                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                    if (_T_443) begin
                                                                                                                                                                                                                                                                                                      bmem_data <= 32'h2c12083;
                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                      if (_T_446) begin
                                                                                                                                                                                                                                                                                                        bmem_data <= 32'h2812403;
                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                        if (_T_449) begin
                                                                                                                                                                                                                                                                                                          bmem_data <= 32'h3010113;
                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                          if (_T_452) begin
                                                                                                                                                                                                                                                                                                            bmem_data <= 32'h8067;
                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                            if (_T_455) begin
                                                                                                                                                                                                                                                                                                              bmem_data <= 32'hfd010113;
                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                              if (_T_458) begin
                                                                                                                                                                                                                                                                                                                bmem_data <= 32'h2112623;
                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                if (_T_461) begin
                                                                                                                                                                                                                                                                                                                  bmem_data <= 32'h2812423;
                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                  if (_T_464) begin
                                                                                                                                                                                                                                                                                                                    bmem_data <= 32'h3010413;
                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                    if (_T_467) begin
                                                                                                                                                                                                                                                                                                                      bmem_data <= 32'hfca42e23;
                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                      if (_T_470) begin
                                                                                                                                                                                                                                                                                                                        bmem_data <= 32'h37b7;
                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                        if (_T_473) begin
                                                                                                                                                                                                                                                                                                                          bmem_data <= 32'h57c783;
                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                          if (_T_476) begin
                                                                                                                                                                                                                                                                                                                            bmem_data <= 32'hff7f713;
                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                            if (_T_479) begin
                                                                                                                                                                                                                                                                                                                              bmem_data <= 32'h37b7;
                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                              if (_T_482) begin
                                                                                                                                                                                                                                                                                                                                bmem_data <= 32'h176713;
                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                if (_T_485) begin
                                                                                                                                                                                                                                                                                                                                  bmem_data <= 32'hff77713;
                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                  if (_T_488) begin
                                                                                                                                                                                                                                                                                                                                    bmem_data <= 32'he782a3;
                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                    if (_T_491) begin
                                                                                                                                                                                                                                                                                                                                      bmem_data <= 32'h300513;
                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                      if (_T_494) begin
                                                                                                                                                                                                                                                                                                                                        bmem_data <= 32'hde1ff0ef;
                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                        if (_T_497) begin
                                                                                                                                                                                                                                                                                                                                          bmem_data <= 32'hfdc42503;
                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                          if (_T_500) begin
                                                                                                                                                                                                                                                                                                                                            bmem_data <= 32'h78000ef;
                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                            if (_T_503) begin
                                                                                                                                                                                                                                                                                                                                              bmem_data <= 32'hfe042623;
                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                              if (_T_506) begin
                                                                                                                                                                                                                                                                                                                                                bmem_data <= 32'h300006f;
                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                if (_T_509) begin
                                                                                                                                                                                                                                                                                                                                                  bmem_data <= 32'h513;
                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                  if (_T_512) begin
                                                                                                                                                                                                                                                                                                                                                    bmem_data <= 32'hdc9ff0ef;
                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                    if (_T_515) begin
                                                                                                                                                                                                                                                                                                                                                      bmem_data <= 32'h50793;
                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                      if (_T_518) begin
                                                                                                                                                                                                                                                                                                                                                        bmem_data <= 32'h78713;
                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                        if (_T_521) begin
                                                                                                                                                                                                                                                                                                                                                          bmem_data <= 32'hfec42783;
                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                          if (_T_524) begin
                                                                                                                                                                                                                                                                                                                                                            bmem_data <= 32'hff040693;
                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                            if (_T_527) begin
                                                                                                                                                                                                                                                                                                                                                              bmem_data <= 32'hf687b3;
                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                              if (_T_530) begin
                                                                                                                                                                                                                                                                                                                                                                bmem_data <= 32'hfee78c23;
                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                if (_T_533) begin
                                                                                                                                                                                                                                                                                                                                                                  bmem_data <= 32'hfec42783;
                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                  if (_T_536) begin
                                                                                                                                                                                                                                                                                                                                                                    bmem_data <= 32'h178793;
                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                    if (_T_539) begin
                                                                                                                                                                                                                                                                                                                                                                      bmem_data <= 32'hfef42623;
                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                      if (_T_542) begin
                                                                                                                                                                                                                                                                                                                                                                        bmem_data <= 32'hfec42703;
                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                        if (_T_545) begin
                                                                                                                                                                                                                                                                                                                                                                          bmem_data <= 32'h300793;
                                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                                          if (_T_548) begin
                                                                                                                                                                                                                                                                                                                                                                            bmem_data <= 32'hfce7f6e3;
                                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                                            if (_T_551) begin
                                                                                                                                                                                                                                                                                                                                                                              bmem_data <= 32'h37b7;
                                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                                              if (_T_554) begin
                                                                                                                                                                                                                                                                                                                                                                                bmem_data <= 32'h57c783;
                                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                                if (_T_557) begin
                                                                                                                                                                                                                                                                                                                                                                                  bmem_data <= 32'hff7f713;
                                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                                  if (_T_560) begin
                                                                                                                                                                                                                                                                                                                                                                                    bmem_data <= 32'h37b7;
                                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                                    if (_T_563) begin
                                                                                                                                                                                                                                                                                                                                                                                      bmem_data <= 32'hffe77713;
                                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                                      if (_T_566) begin
                                                                                                                                                                                                                                                                                                                                                                                        bmem_data <= 32'hff77713;
                                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                                        if (_T_569) begin
                                                                                                                                                                                                                                                                                                                                                                                          bmem_data <= 32'he782a3;
                                                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                                                          if (_T_572) begin
                                                                                                                                                                                                                                                                                                                                                                                            bmem_data <= 32'hfe842783;
                                                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                                                            if (_T_575) begin
                                                                                                                                                                                                                                                                                                                                                                                              bmem_data <= 32'h78513;
                                                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                                                              if (_T_578) begin
                                                                                                                                                                                                                                                                                                                                                                                                bmem_data <= 32'h2c12083;
                                                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                                                if (_T_581) begin
                                                                                                                                                                                                                                                                                                                                                                                                  bmem_data <= 32'h2812403;
                                                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                                                  if (_T_584) begin
                                                                                                                                                                                                                                                                                                                                                                                                    bmem_data <= 32'h3010113;
                                                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                                                    if (_T_587) begin
                                                                                                                                                                                                                                                                                                                                                                                                      bmem_data <= 32'h8067;
                                                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                                                      if (_T_590) begin
                                                                                                                                                                                                                                                                                                                                                                                                        bmem_data <= 32'hfd010113;
                                                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                                                        if (_T_593) begin
                                                                                                                                                                                                                                                                                                                                                                                                          bmem_data <= 32'h2112623;
                                                                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                                                                          if (_T_596) begin
                                                                                                                                                                                                                                                                                                                                                                                                            bmem_data <= 32'h2812423;
                                                                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                                                                            if (_T_599) begin
                                                                                                                                                                                                                                                                                                                                                                                                              bmem_data <= 32'h3010413;
                                                                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                                                                              if (_T_602) begin
                                                                                                                                                                                                                                                                                                                                                                                                                bmem_data <= 32'hfca42e23;
                                                                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                if (_T_605) begin
                                                                                                                                                                                                                                                                                                                                                                                                                  bmem_data <= 32'hfdc42783;
                                                                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                  if (_T_608) begin
                                                                                                                                                                                                                                                                                                                                                                                                                    bmem_data <= 32'hfef42423;
                                                                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                    if (_T_611) begin
                                                                                                                                                                                                                                                                                                                                                                                                                      bmem_data <= 32'h200793;
                                                                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                      if (_T_614) begin
                                                                                                                                                                                                                                                                                                                                                                                                                        bmem_data <= 32'hfef42623;
                                                                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                        if (_T_617) begin
                                                                                                                                                                                                                                                                                                                                                                                                                          bmem_data <= 32'h280006f;
                                                                                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                          if (_T_620) begin
                                                                                                                                                                                                                                                                                                                                                                                                                            bmem_data <= 32'hfec42783;
                                                                                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                            if (_T_623) begin
                                                                                                                                                                                                                                                                                                                                                                                                                              bmem_data <= 32'hff040713;
                                                                                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                              if (_T_626) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                bmem_data <= 32'hf707b3;
                                                                                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                if (_T_629) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                  bmem_data <= 32'hff87c783;
                                                                                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                  if (_T_632) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                    bmem_data <= 32'h78513;
                                                                                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                    if (_T_635) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                      bmem_data <= 32'hd25ff0ef;
                                                                                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                      if (_T_638) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                        bmem_data <= 32'hfec42783;
                                                                                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                        if (_T_641) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                          bmem_data <= 32'hfff78793;
                                                                                                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                          if (_T_644) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                            bmem_data <= 32'hfef42623;
                                                                                                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                            if (_T_647) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                              bmem_data <= 32'hfec42783;
                                                                                                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                              if (_T_650) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                bmem_data <= 32'hfc07dce3;
                                                                                                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                if (_T_653) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                  bmem_data <= 32'h13;
                                                                                                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                  if (_T_656) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                    bmem_data <= 32'h2c12083;
                                                                                                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                    if (_T_659) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                      bmem_data <= 32'h2812403;
                                                                                                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                      if (_T_662) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                        bmem_data <= 32'h3010113;
                                                                                                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                        if (_T_665) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                          bmem_data <= 32'h8067;
                                                                                                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                              end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                          end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                      end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                  end
                                                                                                                                                                                                                end
                                                                                                                                                                                                              end
                                                                                                                                                                                                            end
                                                                                                                                                                                                          end
                                                                                                                                                                                                        end
                                                                                                                                                                                                      end
                                                                                                                                                                                                    end
                                                                                                                                                                                                  end
                                                                                                                                                                                                end
                                                                                                                                                                                              end
                                                                                                                                                                                            end
                                                                                                                                                                                          end
                                                                                                                                                                                        end
                                                                                                                                                                                      end
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end
                                                                                                                                                      end
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end
                                                                                                                                        end
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
