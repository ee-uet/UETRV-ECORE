magic
tech sky130A
magscale 1 2
timestamp 1647908327
<< metal1 >>
rect 204254 325660 204260 325712
rect 204312 325700 204318 325712
rect 207014 325700 207020 325712
rect 204312 325672 207020 325700
rect 204312 325660 204318 325672
rect 207014 325660 207020 325672
rect 207072 325660 207078 325712
rect 193214 306348 193220 306400
rect 193272 306388 193278 306400
rect 207014 306388 207020 306400
rect 193272 306360 207020 306388
rect 193272 306348 193278 306360
rect 207014 306348 207020 306360
rect 207072 306348 207078 306400
rect 190454 304988 190460 305040
rect 190512 305028 190518 305040
rect 207014 305028 207020 305040
rect 190512 305000 207020 305028
rect 190512 304988 190518 305000
rect 207014 304988 207020 305000
rect 207072 304988 207078 305040
rect 55214 298120 55220 298172
rect 55272 298160 55278 298172
rect 55858 298160 55864 298172
rect 55272 298132 55864 298160
rect 55272 298120 55278 298132
rect 55858 298120 55864 298132
rect 55916 298160 55922 298172
rect 215846 298160 215852 298172
rect 55916 298132 215852 298160
rect 55916 298120 55922 298132
rect 215846 298120 215852 298132
rect 215904 298120 215910 298172
rect 95142 297508 95148 297560
rect 95200 297548 95206 297560
rect 130378 297548 130384 297560
rect 95200 297520 130384 297548
rect 95200 297508 95206 297520
rect 130378 297508 130384 297520
rect 130436 297508 130442 297560
rect 71498 297440 71504 297492
rect 71556 297480 71562 297492
rect 130470 297480 130476 297492
rect 71556 297452 130476 297480
rect 71556 297440 71562 297452
rect 130470 297440 130476 297452
rect 130528 297440 130534 297492
rect 81802 297372 81808 297424
rect 81860 297412 81866 297424
rect 188522 297412 188528 297424
rect 81860 297384 188528 297412
rect 81860 297372 81866 297384
rect 188522 297372 188528 297384
rect 188580 297372 188586 297424
rect 76834 297304 76840 297356
rect 76892 297344 76898 297356
rect 188430 297344 188436 297356
rect 76892 297316 188436 297344
rect 76892 297304 76898 297316
rect 188430 297304 188436 297316
rect 188488 297304 188494 297356
rect 65702 297236 65708 297288
rect 65760 297276 65766 297288
rect 188338 297276 188344 297288
rect 65760 297248 188344 297276
rect 65760 297236 65766 297248
rect 188338 297236 188344 297248
rect 188396 297236 188402 297288
rect 67818 297168 67824 297220
rect 67876 297208 67882 297220
rect 227714 297208 227720 297220
rect 67876 297180 227720 297208
rect 67876 297168 67882 297180
rect 227714 297168 227720 297180
rect 227772 297168 227778 297220
rect 70210 297100 70216 297152
rect 70268 297140 70274 297152
rect 229094 297140 229100 297152
rect 70268 297112 229100 297140
rect 70268 297100 70274 297112
rect 229094 297100 229100 297112
rect 229152 297140 229158 297152
rect 229462 297140 229468 297152
rect 229152 297112 229468 297140
rect 229152 297100 229158 297112
rect 229462 297100 229468 297112
rect 229520 297100 229526 297152
rect 69934 297032 69940 297084
rect 69992 297072 69998 297084
rect 229186 297072 229192 297084
rect 69992 297044 229192 297072
rect 69992 297032 69998 297044
rect 229186 297032 229192 297044
rect 229244 297032 229250 297084
rect 79778 296964 79784 297016
rect 79836 297004 79842 297016
rect 352558 297004 352564 297016
rect 79836 296976 352564 297004
rect 79836 296964 79842 296976
rect 352558 296964 352564 296976
rect 352616 296964 352622 297016
rect 106734 296896 106740 296948
rect 106792 296936 106798 296948
rect 409138 296936 409144 296948
rect 106792 296908 409144 296936
rect 106792 296896 106798 296908
rect 409138 296896 409144 296908
rect 409196 296896 409202 296948
rect 103238 296828 103244 296880
rect 103296 296868 103302 296880
rect 409046 296868 409052 296880
rect 103296 296840 409052 296868
rect 103296 296828 103302 296840
rect 409046 296828 409052 296840
rect 409104 296828 409110 296880
rect 96706 296760 96712 296812
rect 96764 296800 96770 296812
rect 408954 296800 408960 296812
rect 96764 296772 408960 296800
rect 96764 296760 96770 296772
rect 408954 296760 408960 296772
rect 409012 296760 409018 296812
rect 93302 296692 93308 296744
rect 93360 296732 93366 296744
rect 408862 296732 408868 296744
rect 93360 296704 408868 296732
rect 93360 296692 93366 296704
rect 408862 296692 408868 296704
rect 408920 296692 408926 296744
rect 267458 263236 267464 263288
rect 267516 263276 267522 263288
rect 371326 263276 371332 263288
rect 267516 263248 371332 263276
rect 267516 263236 267522 263248
rect 371326 263236 371332 263248
rect 371384 263236 371390 263288
rect 110322 263168 110328 263220
rect 110380 263208 110386 263220
rect 411622 263208 411628 263220
rect 110380 263180 411628 263208
rect 110380 263168 110386 263180
rect 411622 263168 411628 263180
rect 411680 263168 411686 263220
rect 104710 263100 104716 263152
rect 104768 263140 104774 263152
rect 410426 263140 410432 263152
rect 104768 263112 410432 263140
rect 104768 263100 104774 263112
rect 410426 263100 410432 263112
rect 410484 263100 410490 263152
rect 99190 263032 99196 263084
rect 99248 263072 99254 263084
rect 411530 263072 411536 263084
rect 99248 263044 411536 263072
rect 99248 263032 99254 263044
rect 411530 263032 411536 263044
rect 411588 263032 411594 263084
rect 86678 262964 86684 263016
rect 86736 263004 86742 263016
rect 409966 263004 409972 263016
rect 86736 262976 409972 263004
rect 86736 262964 86742 262976
rect 409966 262964 409972 262976
rect 410024 262964 410030 263016
rect 81250 262896 81256 262948
rect 81308 262936 81314 262948
rect 410058 262936 410064 262948
rect 81308 262908 410064 262936
rect 81308 262896 81314 262908
rect 410058 262896 410064 262908
rect 410116 262896 410122 262948
rect 75822 262828 75828 262880
rect 75880 262868 75886 262880
rect 411714 262868 411720 262880
rect 75880 262840 411720 262868
rect 75880 262828 75886 262840
rect 411714 262828 411720 262840
rect 411772 262828 411778 262880
rect 259178 261876 259184 261928
rect 259236 261916 259242 261928
rect 338114 261916 338120 261928
rect 259236 261888 338120 261916
rect 259236 261876 259242 261888
rect 338114 261876 338120 261888
rect 338172 261876 338178 261928
rect 263410 261808 263416 261860
rect 263468 261848 263474 261860
rect 352098 261848 352104 261860
rect 263468 261820 352104 261848
rect 263468 261808 263474 261820
rect 352098 261808 352104 261820
rect 352156 261808 352162 261860
rect 264790 261740 264796 261792
rect 264848 261780 264854 261792
rect 356698 261780 356704 261792
rect 264848 261752 356704 261780
rect 264848 261740 264854 261752
rect 356698 261740 356704 261752
rect 356756 261740 356762 261792
rect 266170 261672 266176 261724
rect 266228 261712 266234 261724
rect 361574 261712 361580 261724
rect 266228 261684 361580 261712
rect 266228 261672 266234 261684
rect 361574 261672 361580 261684
rect 361632 261672 361638 261724
rect 267550 261604 267556 261656
rect 267608 261644 267614 261656
rect 366082 261644 366088 261656
rect 267608 261616 366088 261644
rect 267608 261604 267614 261616
rect 366082 261604 366088 261616
rect 366140 261604 366146 261656
rect 104802 261536 104808 261588
rect 104860 261576 104866 261588
rect 406010 261576 406016 261588
rect 104860 261548 406016 261576
rect 104860 261536 104866 261548
rect 406010 261536 406016 261548
rect 406068 261536 406074 261588
rect 81342 261468 81348 261520
rect 81400 261508 81406 261520
rect 385034 261508 385040 261520
rect 81400 261480 385040 261508
rect 81400 261468 81406 261480
rect 385034 261468 385040 261480
rect 385092 261468 385098 261520
rect 253750 260584 253756 260636
rect 253808 260624 253814 260636
rect 314746 260624 314752 260636
rect 253808 260596 314752 260624
rect 253808 260584 253814 260596
rect 314746 260584 314752 260596
rect 314804 260584 314810 260636
rect 255130 260516 255136 260568
rect 255188 260556 255194 260568
rect 319346 260556 319352 260568
rect 255188 260528 319352 260556
rect 255188 260516 255194 260528
rect 319346 260516 319352 260528
rect 319404 260516 319410 260568
rect 256510 260448 256516 260500
rect 256568 260488 256574 260500
rect 324314 260488 324320 260500
rect 256568 260460 324320 260488
rect 256568 260448 256574 260460
rect 324314 260448 324320 260460
rect 324372 260448 324378 260500
rect 257798 260380 257804 260432
rect 257856 260420 257862 260432
rect 328730 260420 328736 260432
rect 257856 260392 328736 260420
rect 257856 260380 257862 260392
rect 328730 260380 328736 260392
rect 328788 260380 328794 260432
rect 259270 260312 259276 260364
rect 259328 260352 259334 260364
rect 333330 260352 333336 260364
rect 259328 260324 333336 260352
rect 259328 260312 259334 260324
rect 333330 260312 333336 260324
rect 333388 260312 333394 260364
rect 260650 260244 260656 260296
rect 260708 260284 260714 260296
rect 342714 260284 342720 260296
rect 260708 260256 342720 260284
rect 260708 260244 260714 260256
rect 342714 260244 342720 260256
rect 342772 260244 342778 260296
rect 79870 260176 79876 260228
rect 79928 260216 79934 260228
rect 378134 260216 378140 260228
rect 79928 260188 378140 260216
rect 79928 260176 79934 260188
rect 378134 260176 378140 260188
rect 378192 260176 378198 260228
rect 100570 260108 100576 260160
rect 100628 260148 100634 260160
rect 401594 260148 401600 260160
rect 100628 260120 401600 260148
rect 100628 260108 100634 260120
rect 401594 260108 401600 260120
rect 401652 260108 401658 260160
rect 246758 259020 246764 259072
rect 246816 259060 246822 259072
rect 286594 259060 286600 259072
rect 246816 259032 286600 259060
rect 246816 259020 246822 259032
rect 286594 259020 286600 259032
rect 286652 259020 286658 259072
rect 248230 258952 248236 259004
rect 248288 258992 248294 259004
rect 291194 258992 291200 259004
rect 248288 258964 291200 258992
rect 248288 258952 248294 258964
rect 291194 258952 291200 258964
rect 291252 258952 291258 259004
rect 249610 258884 249616 258936
rect 249668 258924 249674 258936
rect 295978 258924 295984 258936
rect 249668 258896 295984 258924
rect 249668 258884 249674 258896
rect 295978 258884 295984 258896
rect 296036 258884 296042 258936
rect 250990 258816 250996 258868
rect 251048 258856 251054 258868
rect 300854 258856 300860 258868
rect 251048 258828 300860 258856
rect 251048 258816 251054 258828
rect 300854 258816 300860 258828
rect 300912 258816 300918 258868
rect 252278 258748 252284 258800
rect 252336 258788 252342 258800
rect 305362 258788 305368 258800
rect 252336 258760 305368 258788
rect 252336 258748 252342 258760
rect 305362 258748 305368 258760
rect 305420 258748 305426 258800
rect 262030 258680 262036 258732
rect 262088 258720 262094 258732
rect 347774 258720 347780 258732
rect 262088 258692 347780 258720
rect 262088 258680 262094 258692
rect 347774 258680 347780 258692
rect 347832 258680 347838 258732
rect 245562 257796 245568 257848
rect 245620 257836 245626 257848
rect 282086 257836 282092 257848
rect 245620 257808 282092 257836
rect 245620 257796 245626 257808
rect 282086 257796 282092 257808
rect 282144 257796 282150 257848
rect 260742 257728 260748 257780
rect 260800 257768 260806 257780
rect 307754 257768 307760 257780
rect 260800 257740 307760 257768
rect 260800 257728 260806 257740
rect 307754 257728 307760 257740
rect 307812 257728 307818 257780
rect 262122 257660 262128 257712
rect 262180 257700 262186 257712
rect 312446 257700 312452 257712
rect 262180 257672 312452 257700
rect 262180 257660 262186 257672
rect 312446 257660 312452 257672
rect 312504 257660 312510 257712
rect 263502 257592 263508 257644
rect 263560 257632 263566 257644
rect 317506 257632 317512 257644
rect 263560 257604 317512 257632
rect 263560 257592 263566 257604
rect 317506 257592 317512 257604
rect 317564 257592 317570 257644
rect 266262 257524 266268 257576
rect 266320 257564 266326 257576
rect 326430 257564 326436 257576
rect 266320 257536 326436 257564
rect 266320 257524 266326 257536
rect 326430 257524 326436 257536
rect 326488 257524 326494 257576
rect 273070 257456 273076 257508
rect 273128 257496 273134 257508
rect 354766 257496 354772 257508
rect 273128 257468 354772 257496
rect 273128 257456 273134 257468
rect 354766 257456 354772 257468
rect 354824 257456 354830 257508
rect 90910 257388 90916 257440
rect 90968 257428 90974 257440
rect 410334 257428 410340 257440
rect 90968 257400 410340 257428
rect 90968 257388 90974 257400
rect 410334 257388 410340 257400
rect 410392 257388 410398 257440
rect 78490 257320 78496 257372
rect 78548 257360 78554 257372
rect 409874 257360 409880 257372
rect 78548 257332 409880 257360
rect 78548 257320 78554 257332
rect 409874 257320 409880 257332
rect 409932 257320 409938 257372
rect 242802 256504 242808 256556
rect 242860 256544 242866 256556
rect 268010 256544 268016 256556
rect 242860 256516 268016 256544
rect 242860 256504 242866 256516
rect 268010 256504 268016 256516
rect 268068 256504 268074 256556
rect 255222 256436 255228 256488
rect 255280 256476 255286 256488
rect 284294 256476 284300 256488
rect 255280 256448 284300 256476
rect 255280 256436 255286 256448
rect 284294 256436 284300 256448
rect 284352 256436 284358 256488
rect 219250 256368 219256 256420
rect 219308 256408 219314 256420
rect 229186 256408 229192 256420
rect 219308 256380 229192 256408
rect 219308 256368 219314 256380
rect 229186 256368 229192 256380
rect 229244 256368 229250 256420
rect 256602 256368 256608 256420
rect 256660 256408 256666 256420
rect 289078 256408 289084 256420
rect 256660 256380 289084 256408
rect 256660 256368 256666 256380
rect 289078 256368 289084 256380
rect 289136 256368 289142 256420
rect 210050 256300 210056 256352
rect 210108 256340 210114 256352
rect 227714 256340 227720 256352
rect 210108 256312 227720 256340
rect 210108 256300 210114 256312
rect 227714 256300 227720 256312
rect 227772 256300 227778 256352
rect 257890 256300 257896 256352
rect 257948 256340 257954 256352
rect 293954 256340 293960 256352
rect 257948 256312 293960 256340
rect 257948 256300 257954 256312
rect 293954 256300 293960 256312
rect 294012 256300 294018 256352
rect 212442 256232 212448 256284
rect 212500 256272 212506 256284
rect 231854 256272 231860 256284
rect 212500 256244 231860 256272
rect 212500 256232 212506 256244
rect 231854 256232 231860 256244
rect 231912 256232 231918 256284
rect 257982 256232 257988 256284
rect 258040 256272 258046 256284
rect 298462 256272 298468 256284
rect 258040 256244 298468 256272
rect 258040 256232 258046 256244
rect 298462 256232 298468 256244
rect 298520 256232 298526 256284
rect 201402 256164 201408 256216
rect 201460 256204 201466 256216
rect 226334 256204 226340 256216
rect 201460 256176 226340 256204
rect 201460 256164 201466 256176
rect 226334 256164 226340 256176
rect 226392 256164 226398 256216
rect 259362 256164 259368 256216
rect 259420 256204 259426 256216
rect 303062 256204 303068 256216
rect 259420 256176 303068 256204
rect 259420 256164 259426 256176
rect 303062 256164 303068 256176
rect 303120 256164 303126 256216
rect 93670 256096 93676 256148
rect 93728 256136 93734 256148
rect 250346 256136 250352 256148
rect 93728 256108 250352 256136
rect 93728 256096 93734 256108
rect 250346 256096 250352 256108
rect 250404 256096 250410 256148
rect 277302 256096 277308 256148
rect 277360 256136 277366 256148
rect 368566 256136 368572 256148
rect 277360 256108 368572 256136
rect 277360 256096 277366 256108
rect 368566 256096 368572 256108
rect 368624 256096 368630 256148
rect 49602 256028 49608 256080
rect 49660 256068 49666 256080
rect 387334 256068 387340 256080
rect 49660 256040 387340 256068
rect 49660 256028 49666 256040
rect 387334 256028 387340 256040
rect 387392 256028 387398 256080
rect 47946 255960 47952 256012
rect 48004 256000 48010 256012
rect 410242 256000 410248 256012
rect 48004 255972 410248 256000
rect 48004 255960 48010 255972
rect 410242 255960 410248 255972
rect 410300 255960 410306 256012
rect 217042 255008 217048 255060
rect 217100 255048 217106 255060
rect 240134 255048 240140 255060
rect 217100 255020 240140 255048
rect 217100 255008 217106 255020
rect 240134 255008 240140 255020
rect 240192 255008 240198 255060
rect 252462 255008 252468 255060
rect 252520 255048 252526 255060
rect 274910 255048 274916 255060
rect 252520 255020 274916 255048
rect 252520 255008 252526 255020
rect 274910 255008 274916 255020
rect 274968 255008 274974 255060
rect 202690 254940 202696 254992
rect 202748 254980 202754 254992
rect 230474 254980 230480 254992
rect 202748 254952 230480 254980
rect 202748 254940 202754 254952
rect 230474 254940 230480 254952
rect 230532 254940 230538 254992
rect 253842 254940 253848 254992
rect 253900 254980 253906 254992
rect 279694 254980 279700 254992
rect 253900 254952 279700 254980
rect 253900 254940 253906 254952
rect 279694 254940 279700 254952
rect 279752 254940 279758 254992
rect 209590 254872 209596 254924
rect 209648 254912 209654 254924
rect 240134 254912 240140 254924
rect 209648 254884 240140 254912
rect 209648 254872 209654 254884
rect 240134 254872 240140 254884
rect 240192 254872 240198 254924
rect 244090 254872 244096 254924
rect 244148 254912 244154 254924
rect 277486 254912 277492 254924
rect 244148 254884 277492 254912
rect 244148 254872 244154 254884
rect 277486 254872 277492 254884
rect 277544 254872 277550 254924
rect 207842 254804 207848 254856
rect 207900 254844 207906 254856
rect 238754 254844 238760 254856
rect 207900 254816 238760 254844
rect 207900 254804 207906 254816
rect 238754 254804 238760 254816
rect 238812 254804 238818 254856
rect 252370 254804 252376 254856
rect 252428 254844 252434 254856
rect 310054 254844 310060 254856
rect 252428 254816 310060 254844
rect 252428 254804 252434 254816
rect 310054 254804 310060 254816
rect 310112 254804 310118 254856
rect 209682 254736 209688 254788
rect 209740 254776 209746 254788
rect 247034 254776 247040 254788
rect 209740 254748 247040 254776
rect 209740 254736 209746 254748
rect 247034 254736 247040 254748
rect 247092 254736 247098 254788
rect 251082 254736 251088 254788
rect 251140 254776 251146 254788
rect 270494 254776 270500 254788
rect 251140 254748 270500 254776
rect 251140 254736 251146 254748
rect 270494 254736 270500 254748
rect 270552 254736 270558 254788
rect 273162 254736 273168 254788
rect 273220 254776 273226 254788
rect 349798 254776 349804 254788
rect 273220 254748 349804 254776
rect 273220 254736 273226 254748
rect 349798 254736 349804 254748
rect 349856 254736 349862 254788
rect 47670 254668 47676 254720
rect 47728 254708 47734 254720
rect 373350 254708 373356 254720
rect 47728 254680 373356 254708
rect 47728 254668 47734 254680
rect 373350 254668 373356 254680
rect 373408 254668 373414 254720
rect 47762 254600 47768 254652
rect 47820 254640 47826 254652
rect 382550 254640 382556 254652
rect 47820 254612 382556 254640
rect 47820 254600 47826 254612
rect 382550 254600 382556 254612
rect 382608 254600 382614 254652
rect 47854 254532 47860 254584
rect 47912 254572 47918 254584
rect 410150 254572 410156 254584
rect 47912 254544 410156 254572
rect 47912 254532 47918 254544
rect 410150 254532 410156 254544
rect 410208 254532 410214 254584
rect 228726 253852 228732 253904
rect 228784 253892 228790 253904
rect 229094 253892 229100 253904
rect 228784 253864 229100 253892
rect 228784 253852 228790 253864
rect 229094 253852 229100 253864
rect 229152 253852 229158 253904
rect 246942 253852 246948 253904
rect 247000 253892 247006 253904
rect 249150 253892 249156 253904
rect 247000 253864 249156 253892
rect 247000 253852 247006 253864
rect 249150 253852 249156 253864
rect 249208 253852 249214 253904
rect 242802 253784 242808 253836
rect 242860 253824 242866 253836
rect 244274 253824 244280 253836
rect 242860 253796 244280 253824
rect 242860 253784 242866 253796
rect 244274 253784 244280 253796
rect 244332 253784 244338 253836
rect 264882 253580 264888 253632
rect 264940 253620 264946 253632
rect 321830 253620 321836 253632
rect 264940 253592 321836 253620
rect 264940 253580 264946 253592
rect 321830 253580 321836 253592
rect 321888 253580 321894 253632
rect 208026 253512 208032 253564
rect 208084 253552 208090 253564
rect 214190 253552 214196 253564
rect 208084 253524 214196 253552
rect 208084 253512 208090 253524
rect 214190 253512 214196 253524
rect 214248 253512 214254 253564
rect 221826 253512 221832 253564
rect 221884 253552 221890 253564
rect 233234 253552 233240 253564
rect 221884 253524 233240 253552
rect 221884 253512 221890 253524
rect 233234 253512 233240 253524
rect 233292 253512 233298 253564
rect 237190 253512 237196 253564
rect 237248 253552 237254 253564
rect 244550 253552 244556 253564
rect 237248 253524 244556 253552
rect 237248 253512 237254 253524
rect 244550 253512 244556 253524
rect 244608 253512 244614 253564
rect 246850 253512 246856 253564
rect 246908 253552 246914 253564
rect 256326 253552 256332 253564
rect 246908 253524 256332 253552
rect 246908 253512 246914 253524
rect 256326 253512 256332 253524
rect 256384 253512 256390 253564
rect 267642 253512 267648 253564
rect 267700 253552 267706 253564
rect 331214 253552 331220 253564
rect 267700 253524 331220 253552
rect 267700 253512 267706 253524
rect 331214 253512 331220 253524
rect 331272 253512 331278 253564
rect 208118 253444 208124 253496
rect 208176 253484 208182 253496
rect 223574 253484 223580 253496
rect 208176 253456 223580 253484
rect 208176 253444 208182 253456
rect 223574 253444 223580 253456
rect 223632 253444 223638 253496
rect 226242 253444 226248 253496
rect 226300 253484 226306 253496
rect 241514 253484 241520 253496
rect 226300 253456 241520 253484
rect 226300 253444 226306 253456
rect 241514 253444 241520 253456
rect 241572 253444 241578 253496
rect 248322 253444 248328 253496
rect 248380 253484 248386 253496
rect 260926 253484 260932 253496
rect 248380 253456 260932 253484
rect 248380 253444 248386 253456
rect 260926 253444 260932 253456
rect 260984 253444 260990 253496
rect 269022 253444 269028 253496
rect 269080 253484 269086 253496
rect 335814 253484 335820 253496
rect 269080 253456 335820 253484
rect 269080 253444 269086 253456
rect 335814 253444 335820 253456
rect 335872 253444 335878 253496
rect 208210 253376 208216 253428
rect 208268 253416 208274 253428
rect 232774 253416 232780 253428
rect 208268 253388 232780 253416
rect 208268 253376 208274 253388
rect 232774 253376 232780 253388
rect 232832 253376 232838 253428
rect 235810 253376 235816 253428
rect 235868 253416 235874 253428
rect 242894 253416 242900 253428
rect 235868 253388 242900 253416
rect 235868 253376 235874 253388
rect 242894 253376 242900 253388
rect 242952 253376 242958 253428
rect 249702 253376 249708 253428
rect 249760 253416 249766 253428
rect 265526 253416 265532 253428
rect 249760 253388 265532 253416
rect 249760 253376 249766 253388
rect 265526 253376 265532 253388
rect 265584 253376 265590 253428
rect 270402 253376 270408 253428
rect 270460 253416 270466 253428
rect 340414 253416 340420 253428
rect 270460 253388 340420 253416
rect 270460 253376 270466 253388
rect 340414 253376 340420 253388
rect 340472 253376 340478 253428
rect 195790 253308 195796 253360
rect 195848 253348 195854 253360
rect 224954 253348 224960 253360
rect 195848 253320 224960 253348
rect 195848 253308 195854 253320
rect 224954 253308 224960 253320
rect 225012 253308 225018 253360
rect 240042 253308 240048 253360
rect 240100 253348 240106 253360
rect 258534 253348 258540 253360
rect 240100 253320 258540 253348
rect 240100 253308 240106 253320
rect 258534 253308 258540 253320
rect 258592 253308 258598 253360
rect 271782 253308 271788 253360
rect 271840 253348 271846 253360
rect 345198 253348 345204 253360
rect 271840 253320 345204 253348
rect 271840 253308 271846 253320
rect 345198 253308 345204 253320
rect 345256 253308 345262 253360
rect 198458 253240 198464 253292
rect 198516 253280 198522 253292
rect 237374 253280 237380 253292
rect 198516 253252 237380 253280
rect 198516 253240 198522 253252
rect 237374 253240 237380 253252
rect 237432 253240 237438 253292
rect 244182 253240 244188 253292
rect 244240 253280 244246 253292
rect 272702 253280 272708 253292
rect 244240 253252 272708 253280
rect 244240 253240 244246 253252
rect 272702 253240 272708 253252
rect 272760 253240 272766 253292
rect 274542 253240 274548 253292
rect 274600 253280 274606 253292
rect 359182 253280 359188 253292
rect 274600 253252 359188 253280
rect 274600 253240 274606 253252
rect 359182 253240 359188 253252
rect 359240 253240 359246 253292
rect 77110 253172 77116 253224
rect 77168 253212 77174 253224
rect 147674 253212 147680 253224
rect 77168 253184 147680 253212
rect 77168 253172 77174 253184
rect 147674 253172 147680 253184
rect 147732 253172 147738 253224
rect 208302 253172 208308 253224
rect 208360 253212 208366 253224
rect 253934 253212 253940 253224
rect 208360 253184 253940 253212
rect 208360 253172 208366 253184
rect 253934 253172 253940 253184
rect 253992 253172 253998 253224
rect 275922 253172 275928 253224
rect 275980 253212 275986 253224
rect 363966 253212 363972 253224
rect 275980 253184 363972 253212
rect 275980 253172 275986 253184
rect 363966 253172 363972 253184
rect 364024 253172 364030 253224
rect 231210 253104 231216 253156
rect 231268 253144 231274 253156
rect 234614 253144 234620 253156
rect 231268 253116 234620 253144
rect 231268 253104 231274 253116
rect 234614 253104 234620 253116
rect 234672 253104 234678 253156
rect 67542 252492 67548 252544
rect 67600 252532 67606 252544
rect 200482 252532 200488 252544
rect 67600 252504 200488 252532
rect 67600 252492 67606 252504
rect 200482 252492 200488 252504
rect 200540 252532 200546 252544
rect 201402 252532 201408 252544
rect 200540 252504 201408 252532
rect 200540 252492 200546 252504
rect 201402 252492 201408 252504
rect 201460 252492 201466 252544
rect 238662 252356 238668 252408
rect 238720 252396 238726 252408
rect 251542 252396 251548 252408
rect 238720 252368 251548 252396
rect 238720 252356 238726 252368
rect 251542 252356 251548 252368
rect 251600 252356 251606 252408
rect 241422 252288 241428 252340
rect 241480 252328 241486 252340
rect 263686 252328 263692 252340
rect 241480 252300 263692 252328
rect 241480 252288 241486 252300
rect 263686 252288 263692 252300
rect 263744 252288 263750 252340
rect 352558 252288 352564 252340
rect 352616 252328 352622 252340
rect 394326 252328 394332 252340
rect 352616 252300 394332 252328
rect 352616 252288 352622 252300
rect 394326 252288 394332 252300
rect 394384 252288 394390 252340
rect 250346 252220 250352 252272
rect 250404 252260 250410 252272
rect 403710 252260 403716 252272
rect 250404 252232 403716 252260
rect 250404 252220 250410 252232
rect 403710 252220 403716 252232
rect 403768 252220 403774 252272
rect 147674 252152 147680 252204
rect 147732 252192 147738 252204
rect 391934 252192 391940 252204
rect 147732 252164 391940 252192
rect 147732 252152 147738 252164
rect 391934 252152 391940 252164
rect 391992 252152 391998 252204
rect 111702 252084 111708 252136
rect 111760 252124 111766 252136
rect 408586 252124 408592 252136
rect 111760 252096 408592 252124
rect 111760 252084 111766 252096
rect 408586 252084 408592 252096
rect 408644 252084 408650 252136
rect 84010 252016 84016 252068
rect 84068 252056 84074 252068
rect 389726 252056 389732 252068
rect 84068 252028 389732 252056
rect 84068 252016 84074 252028
rect 389726 252016 389732 252028
rect 389784 252016 389790 252068
rect 91002 251948 91008 252000
rect 91060 251988 91066 252000
rect 398926 251988 398932 252000
rect 91060 251960 398932 251988
rect 91060 251948 91066 251960
rect 398926 251948 398932 251960
rect 398984 251948 398990 252000
rect 88150 251880 88156 251932
rect 88208 251920 88214 251932
rect 396718 251920 396724 251932
rect 88208 251892 396724 251920
rect 88208 251880 88214 251892
rect 396718 251880 396724 251892
rect 396776 251880 396782 251932
rect 49510 251812 49516 251864
rect 49568 251852 49574 251864
rect 375558 251852 375564 251864
rect 49568 251824 375564 251852
rect 49568 251812 49574 251824
rect 375558 251812 375564 251824
rect 375616 251812 375622 251864
rect 117222 250792 117228 250844
rect 117280 250832 117286 250844
rect 408494 250832 408500 250844
rect 117280 250804 408500 250832
rect 117280 250792 117286 250804
rect 408494 250792 408500 250804
rect 408552 250792 408558 250844
rect 114462 250724 114468 250776
rect 114520 250764 114526 250776
rect 410518 250764 410524 250776
rect 114520 250736 410524 250764
rect 114520 250724 114526 250736
rect 410518 250724 410524 250736
rect 410576 250724 410582 250776
rect 115842 250656 115848 250708
rect 115900 250696 115906 250708
rect 411254 250696 411260 250708
rect 115900 250668 411260 250696
rect 115900 250656 115906 250668
rect 411254 250656 411260 250668
rect 411312 250656 411318 250708
rect 107470 250588 107476 250640
rect 107528 250628 107534 250640
rect 411438 250628 411444 250640
rect 107528 250600 411444 250628
rect 107528 250588 107534 250600
rect 411438 250588 411444 250600
rect 411496 250588 411502 250640
rect 73062 250520 73068 250572
rect 73120 250560 73126 250572
rect 411806 250560 411812 250572
rect 73120 250532 411812 250560
rect 73120 250520 73126 250532
rect 411806 250520 411812 250532
rect 411864 250520 411870 250572
rect 48038 250452 48044 250504
rect 48096 250492 48102 250504
rect 411346 250492 411352 250504
rect 48096 250464 411352 250492
rect 48096 250452 48102 250464
rect 411346 250452 411352 250464
rect 411404 250452 411410 250504
rect 187234 249772 187240 249824
rect 187292 249812 187298 249824
rect 580350 249812 580356 249824
rect 187292 249784 580356 249812
rect 187292 249772 187298 249784
rect 580350 249772 580356 249784
rect 580408 249772 580414 249824
rect 106090 249704 106096 249756
rect 106148 249744 106154 249756
rect 187510 249744 187516 249756
rect 106148 249716 187516 249744
rect 106148 249704 106154 249716
rect 187510 249704 187516 249716
rect 187568 249704 187574 249756
rect 108850 249636 108856 249688
rect 108908 249676 108914 249688
rect 187602 249676 187608 249688
rect 108908 249648 187608 249676
rect 108908 249636 108914 249648
rect 187602 249636 187608 249648
rect 187660 249636 187666 249688
rect 187418 248412 187424 248464
rect 187476 248452 187482 248464
rect 580258 248452 580264 248464
rect 187476 248424 580264 248452
rect 187476 248412 187482 248424
rect 580258 248412 580264 248424
rect 580316 248412 580322 248464
rect 112990 248344 112996 248396
rect 113048 248384 113054 248396
rect 187602 248384 187608 248396
rect 113048 248356 187608 248384
rect 113048 248344 113054 248356
rect 187602 248344 187608 248356
rect 187660 248344 187666 248396
rect 113082 246984 113088 247036
rect 113140 247024 113146 247036
rect 187326 247024 187332 247036
rect 113140 246996 187332 247024
rect 113140 246984 113146 246996
rect 187326 246984 187332 246996
rect 187384 246984 187390 247036
rect 101858 245556 101864 245608
rect 101916 245596 101922 245608
rect 187602 245596 187608 245608
rect 101916 245568 187608 245596
rect 101916 245556 101922 245568
rect 187602 245556 187608 245568
rect 187660 245556 187666 245608
rect 101950 244196 101956 244248
rect 102008 244236 102014 244248
rect 186314 244236 186320 244248
rect 102008 244208 186320 244236
rect 102008 244196 102014 244208
rect 186314 244196 186320 244208
rect 186372 244196 186378 244248
rect 411254 243516 411260 243568
rect 411312 243556 411318 243568
rect 411438 243556 411444 243568
rect 411312 243528 411444 243556
rect 411312 243516 411318 243528
rect 411438 243516 411444 243528
rect 411496 243516 411502 243568
rect 411438 243380 411444 243432
rect 411496 243420 411502 243432
rect 411806 243420 411812 243432
rect 411496 243392 411812 243420
rect 411496 243380 411502 243392
rect 411806 243380 411812 243392
rect 411864 243380 411870 243432
rect 102042 242836 102048 242888
rect 102100 242876 102106 242888
rect 186406 242876 186412 242888
rect 102100 242848 186412 242876
rect 102100 242836 102106 242848
rect 186406 242836 186412 242848
rect 186464 242836 186470 242888
rect 106182 242768 106188 242820
rect 106240 242808 106246 242820
rect 186314 242808 186320 242820
rect 106240 242780 186320 242808
rect 106240 242768 106246 242780
rect 186314 242768 186320 242780
rect 186372 242768 186378 242820
rect 93578 241408 93584 241460
rect 93636 241448 93642 241460
rect 186314 241448 186320 241460
rect 93636 241420 186320 241448
rect 93636 241408 93642 241420
rect 186314 241408 186320 241420
rect 186372 241408 186378 241460
rect 99282 240048 99288 240100
rect 99340 240088 99346 240100
rect 186314 240088 186320 240100
rect 99340 240060 186320 240088
rect 99340 240048 99346 240060
rect 186314 240048 186320 240060
rect 186372 240048 186378 240100
rect 89530 238688 89536 238740
rect 89588 238728 89594 238740
rect 186314 238728 186320 238740
rect 89588 238700 186320 238728
rect 89588 238688 89594 238700
rect 186314 238688 186320 238700
rect 186372 238688 186378 238740
rect 86770 237328 86776 237380
rect 86828 237368 86834 237380
rect 186406 237368 186412 237380
rect 86828 237340 186412 237368
rect 86828 237328 86834 237340
rect 186406 237328 186412 237340
rect 186464 237328 186470 237380
rect 96430 237260 96436 237312
rect 96488 237300 96494 237312
rect 186314 237300 186320 237312
rect 96488 237272 186320 237300
rect 96488 237260 96494 237272
rect 186314 237260 186320 237272
rect 186372 237260 186378 237312
rect 95050 235900 95056 235952
rect 95108 235940 95114 235952
rect 186314 235940 186320 235952
rect 95108 235912 186320 235940
rect 95108 235900 95114 235912
rect 186314 235900 186320 235912
rect 186372 235900 186378 235952
rect 89622 234540 89628 234592
rect 89680 234580 89686 234592
rect 186314 234580 186320 234592
rect 89680 234552 186320 234580
rect 89680 234540 89686 234552
rect 186314 234540 186320 234552
rect 186372 234540 186378 234592
rect 78582 233180 78588 233232
rect 78640 233220 78646 233232
rect 186314 233220 186320 233232
rect 78640 233192 186320 233220
rect 78640 233180 78646 233192
rect 186314 233180 186320 233192
rect 186372 233180 186378 233232
rect 463694 231820 463700 231872
rect 463752 231860 463758 231872
rect 579614 231860 579620 231872
rect 463752 231832 579620 231860
rect 463752 231820 463758 231832
rect 579614 231820 579620 231832
rect 579672 231820 579678 231872
rect 48130 231752 48136 231804
rect 48188 231792 48194 231804
rect 186314 231792 186320 231804
rect 48188 231764 186320 231792
rect 48188 231752 48194 231764
rect 186314 231752 186320 231764
rect 186372 231752 186378 231804
rect 82630 230392 82636 230444
rect 82688 230432 82694 230444
rect 186314 230432 186320 230444
rect 82688 230404 186320 230432
rect 82688 230392 82694 230404
rect 186314 230392 186320 230404
rect 186372 230392 186378 230444
rect 74442 229032 74448 229084
rect 74500 229072 74506 229084
rect 186314 229072 186320 229084
rect 74500 229044 186320 229072
rect 74500 229032 74506 229044
rect 186314 229032 186320 229044
rect 186372 229032 186378 229084
rect 169018 222164 169024 222216
rect 169076 222204 169082 222216
rect 186314 222204 186320 222216
rect 169076 222176 186320 222204
rect 169076 222164 169082 222176
rect 186314 222164 186320 222176
rect 186372 222164 186378 222216
rect 131850 220804 131856 220856
rect 131908 220844 131914 220856
rect 186314 220844 186320 220856
rect 131908 220816 186320 220844
rect 131908 220804 131914 220816
rect 186314 220804 186320 220816
rect 186372 220804 186378 220856
rect 159358 219444 159364 219496
rect 159416 219484 159422 219496
rect 186314 219484 186320 219496
rect 159416 219456 186320 219484
rect 159416 219444 159422 219456
rect 186314 219444 186320 219456
rect 186372 219444 186378 219496
rect 135990 218016 135996 218068
rect 136048 218056 136054 218068
rect 186314 218056 186320 218068
rect 136048 218028 186320 218056
rect 136048 218016 136054 218028
rect 186314 218016 186320 218028
rect 186372 218016 186378 218068
rect 542998 218016 543004 218068
rect 543056 218056 543062 218068
rect 580166 218056 580172 218068
rect 543056 218028 580172 218056
rect 543056 218016 543062 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 142798 216724 142804 216776
rect 142856 216764 142862 216776
rect 186406 216764 186412 216776
rect 142856 216736 186412 216764
rect 142856 216724 142862 216736
rect 186406 216724 186412 216736
rect 186464 216724 186470 216776
rect 135898 216656 135904 216708
rect 135956 216696 135962 216708
rect 186314 216696 186320 216708
rect 135956 216668 186320 216696
rect 135956 216656 135962 216668
rect 186314 216656 186320 216668
rect 186372 216656 186378 216708
rect 157978 215296 157984 215348
rect 158036 215336 158042 215348
rect 186314 215336 186320 215348
rect 158036 215308 186320 215336
rect 158036 215296 158042 215308
rect 186314 215296 186320 215308
rect 186372 215296 186378 215348
rect 134518 213936 134524 213988
rect 134576 213976 134582 213988
rect 186314 213976 186320 213988
rect 134576 213948 186320 213976
rect 134576 213936 134582 213948
rect 186314 213936 186320 213948
rect 186372 213936 186378 213988
rect 141418 212508 141424 212560
rect 141476 212548 141482 212560
rect 186314 212548 186320 212560
rect 141476 212520 186320 212548
rect 141476 212508 141482 212520
rect 186314 212508 186320 212520
rect 186372 212508 186378 212560
rect 156598 211148 156604 211200
rect 156656 211188 156662 211200
rect 186314 211188 186320 211200
rect 156656 211160 186320 211188
rect 156656 211148 156662 211160
rect 186314 211148 186320 211160
rect 186372 211148 186378 211200
rect 136082 209788 136088 209840
rect 136140 209828 136146 209840
rect 186314 209828 186320 209840
rect 136140 209800 186320 209828
rect 136140 209788 136146 209800
rect 186314 209788 186320 209800
rect 186372 209788 186378 209840
rect 411254 209788 411260 209840
rect 411312 209828 411318 209840
rect 418798 209828 418804 209840
rect 411312 209800 418804 209828
rect 411312 209788 411318 209800
rect 418798 209788 418804 209800
rect 418856 209788 418862 209840
rect 141510 208360 141516 208412
rect 141568 208400 141574 208412
rect 186314 208400 186320 208412
rect 141568 208372 186320 208400
rect 141568 208360 141574 208372
rect 186314 208360 186320 208372
rect 186372 208360 186378 208412
rect 133230 207000 133236 207052
rect 133288 207040 133294 207052
rect 186314 207040 186320 207052
rect 133288 207012 186320 207040
rect 133288 207000 133294 207012
rect 186314 207000 186320 207012
rect 186372 207000 186378 207052
rect 411254 207000 411260 207052
rect 411312 207040 411318 207052
rect 414658 207040 414664 207052
rect 411312 207012 414664 207040
rect 411312 207000 411318 207012
rect 414658 207000 414664 207012
rect 414716 207000 414722 207052
rect 155218 205640 155224 205692
rect 155276 205680 155282 205692
rect 186314 205680 186320 205692
rect 155276 205652 186320 205680
rect 155276 205640 155282 205652
rect 186314 205640 186320 205652
rect 186372 205640 186378 205692
rect 411254 205640 411260 205692
rect 411312 205680 411318 205692
rect 544378 205680 544384 205692
rect 411312 205652 544384 205680
rect 411312 205640 411318 205652
rect 544378 205640 544384 205652
rect 544436 205640 544442 205692
rect 142890 204280 142896 204332
rect 142948 204320 142954 204332
rect 186314 204320 186320 204332
rect 142948 204292 186320 204320
rect 142948 204280 142954 204292
rect 186314 204280 186320 204292
rect 186372 204280 186378 204332
rect 134610 202852 134616 202904
rect 134668 202892 134674 202904
rect 186314 202892 186320 202904
rect 134668 202864 186320 202892
rect 134668 202852 134674 202864
rect 186314 202852 186320 202864
rect 186372 202852 186378 202904
rect 411254 202852 411260 202904
rect 411312 202892 411318 202904
rect 540238 202892 540244 202904
rect 411312 202864 540244 202892
rect 411312 202852 411318 202864
rect 540238 202852 540244 202864
rect 540296 202852 540302 202904
rect 152458 201492 152464 201544
rect 152516 201532 152522 201544
rect 186314 201532 186320 201544
rect 152516 201504 186320 201532
rect 152516 201492 152522 201504
rect 186314 201492 186320 201504
rect 186372 201492 186378 201544
rect 134702 200132 134708 200184
rect 134760 200172 134766 200184
rect 186314 200172 186320 200184
rect 134760 200144 186320 200172
rect 134760 200132 134766 200144
rect 186314 200132 186320 200144
rect 186372 200132 186378 200184
rect 151078 198772 151084 198824
rect 151136 198812 151142 198824
rect 186406 198812 186412 198824
rect 151136 198784 186412 198812
rect 151136 198772 151142 198784
rect 186406 198772 186412 198784
rect 186464 198772 186470 198824
rect 134794 198704 134800 198756
rect 134852 198744 134858 198756
rect 186314 198744 186320 198756
rect 134852 198716 186320 198744
rect 134852 198704 134858 198716
rect 186314 198704 186320 198716
rect 186372 198704 186378 198756
rect 148318 197344 148324 197396
rect 148376 197384 148382 197396
rect 186314 197384 186320 197396
rect 148376 197356 186320 197384
rect 148376 197344 148382 197356
rect 186314 197344 186320 197356
rect 186372 197344 186378 197396
rect 411254 197344 411260 197396
rect 411312 197384 411318 197396
rect 421558 197384 421564 197396
rect 411312 197356 421564 197384
rect 411312 197344 411318 197356
rect 421558 197344 421564 197356
rect 421616 197344 421622 197396
rect 134886 195984 134892 196036
rect 134944 196024 134950 196036
rect 186314 196024 186320 196036
rect 134944 195996 186320 196024
rect 134944 195984 134950 195996
rect 186314 195984 186320 195996
rect 186372 195984 186378 196036
rect 411254 195984 411260 196036
rect 411312 196024 411318 196036
rect 416038 196024 416044 196036
rect 411312 195996 416044 196024
rect 411312 195984 411318 195996
rect 416038 195984 416044 195996
rect 416096 195984 416102 196036
rect 145558 194556 145564 194608
rect 145616 194596 145622 194608
rect 186314 194596 186320 194608
rect 145616 194568 186320 194596
rect 145616 194556 145622 194568
rect 186314 194556 186320 194568
rect 186372 194556 186378 194608
rect 134978 193196 134984 193248
rect 135036 193236 135042 193248
rect 186314 193236 186320 193248
rect 135036 193208 186320 193236
rect 135036 193196 135042 193208
rect 186314 193196 186320 193208
rect 186372 193196 186378 193248
rect 146938 191904 146944 191956
rect 146996 191944 147002 191956
rect 186406 191944 186412 191956
rect 146996 191916 186412 191944
rect 146996 191904 147002 191916
rect 186406 191904 186412 191916
rect 186464 191904 186470 191956
rect 133322 191836 133328 191888
rect 133380 191876 133386 191888
rect 186314 191876 186320 191888
rect 133380 191848 186320 191876
rect 133380 191836 133386 191848
rect 186314 191836 186320 191848
rect 186372 191836 186378 191888
rect 411254 191836 411260 191888
rect 411312 191876 411318 191888
rect 436738 191876 436744 191888
rect 411312 191848 436744 191876
rect 411312 191836 411318 191848
rect 436738 191836 436744 191848
rect 436796 191836 436802 191888
rect 543182 191836 543188 191888
rect 543240 191876 543246 191888
rect 580166 191876 580172 191888
rect 543240 191848 580172 191876
rect 543240 191836 543246 191848
rect 580166 191836 580172 191848
rect 580224 191836 580230 191888
rect 147030 190476 147036 190528
rect 147088 190516 147094 190528
rect 186314 190516 186320 190528
rect 147088 190488 186320 190516
rect 147088 190476 147094 190488
rect 186314 190476 186320 190488
rect 186372 190476 186378 190528
rect 145650 189048 145656 189100
rect 145708 189088 145714 189100
rect 186314 189088 186320 189100
rect 145708 189060 186320 189088
rect 145708 189048 145714 189060
rect 186314 189048 186320 189060
rect 186372 189048 186378 189100
rect 411254 189048 411260 189100
rect 411312 189088 411318 189100
rect 421650 189088 421656 189100
rect 411312 189060 421656 189088
rect 411312 189048 411318 189060
rect 421650 189048 421656 189060
rect 421708 189048 421714 189100
rect 140130 187688 140136 187740
rect 140188 187728 140194 187740
rect 186314 187728 186320 187740
rect 140188 187700 186320 187728
rect 140188 187688 140194 187700
rect 186314 187688 186320 187700
rect 186372 187688 186378 187740
rect 411254 187688 411260 187740
rect 411312 187728 411318 187740
rect 435358 187728 435364 187740
rect 411312 187700 435364 187728
rect 411312 187688 411318 187700
rect 435358 187688 435364 187700
rect 435416 187688 435422 187740
rect 140038 186396 140044 186448
rect 140096 186436 140102 186448
rect 186314 186436 186320 186448
rect 140096 186408 186320 186436
rect 140096 186396 140102 186408
rect 186314 186396 186320 186408
rect 186372 186396 186378 186448
rect 133414 186328 133420 186380
rect 133472 186368 133478 186380
rect 186406 186368 186412 186380
rect 133472 186340 186412 186368
rect 133472 186328 133478 186340
rect 186406 186328 186412 186340
rect 186464 186328 186470 186380
rect 411254 184900 411260 184952
rect 411312 184940 411318 184952
rect 416130 184940 416136 184952
rect 411312 184912 416136 184940
rect 411312 184900 411318 184912
rect 416130 184900 416136 184912
rect 416188 184900 416194 184952
rect 137278 183540 137284 183592
rect 137336 183580 137342 183592
rect 186314 183580 186320 183592
rect 137336 183552 186320 183580
rect 137336 183540 137342 183552
rect 186314 183540 186320 183552
rect 186372 183540 186378 183592
rect 411254 183540 411260 183592
rect 411312 183580 411318 183592
rect 432598 183580 432604 183592
rect 411312 183552 432604 183580
rect 411312 183540 411318 183552
rect 432598 183540 432604 183552
rect 432656 183540 432662 183592
rect 145742 182180 145748 182232
rect 145800 182220 145806 182232
rect 186314 182220 186320 182232
rect 145800 182192 186320 182220
rect 145800 182180 145806 182192
rect 186314 182180 186320 182192
rect 186372 182180 186378 182232
rect 411254 182180 411260 182232
rect 411312 182220 411318 182232
rect 431218 182220 431224 182232
rect 411312 182192 431224 182220
rect 411312 182180 411318 182192
rect 431218 182180 431224 182192
rect 431276 182180 431282 182232
rect 140222 180820 140228 180872
rect 140280 180860 140286 180872
rect 186314 180860 186320 180872
rect 140280 180832 186320 180860
rect 140280 180820 140286 180832
rect 186314 180820 186320 180832
rect 186372 180820 186378 180872
rect 140314 179460 140320 179512
rect 140372 179500 140378 179512
rect 186314 179500 186320 179512
rect 140372 179472 186320 179500
rect 140372 179460 140378 179472
rect 186314 179460 186320 179472
rect 186372 179460 186378 179512
rect 133598 179392 133604 179444
rect 133656 179432 133662 179444
rect 186406 179432 186412 179444
rect 133656 179404 186412 179432
rect 133656 179392 133662 179404
rect 186406 179392 186412 179404
rect 186464 179392 186470 179444
rect 411254 179392 411260 179444
rect 411312 179432 411318 179444
rect 429838 179432 429844 179444
rect 411312 179404 429844 179432
rect 411312 179392 411318 179404
rect 429838 179392 429844 179404
rect 429896 179392 429902 179444
rect 133506 178032 133512 178084
rect 133564 178072 133570 178084
rect 186314 178072 186320 178084
rect 133564 178044 186320 178072
rect 133564 178032 133570 178044
rect 186314 178032 186320 178044
rect 186372 178032 186378 178084
rect 411254 178032 411260 178084
rect 411312 178072 411318 178084
rect 428458 178072 428464 178084
rect 411312 178044 428464 178072
rect 411312 178032 411318 178044
rect 428458 178032 428464 178044
rect 428516 178032 428522 178084
rect 543090 178032 543096 178084
rect 543148 178072 543154 178084
rect 580166 178072 580172 178084
rect 543148 178044 580172 178072
rect 543148 178032 543154 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 138658 176672 138664 176724
rect 138716 176712 138722 176724
rect 186314 176712 186320 176724
rect 138716 176684 186320 176712
rect 138716 176672 138722 176684
rect 186314 176672 186320 176684
rect 186372 176672 186378 176724
rect 133690 175244 133696 175296
rect 133748 175284 133754 175296
rect 186314 175284 186320 175296
rect 133748 175256 186320 175284
rect 133748 175244 133754 175256
rect 186314 175244 186320 175256
rect 186372 175244 186378 175296
rect 411254 175244 411260 175296
rect 411312 175284 411318 175296
rect 425698 175284 425704 175296
rect 411312 175256 425704 175284
rect 411312 175244 411318 175256
rect 425698 175244 425704 175256
rect 425756 175244 425762 175296
rect 137370 173884 137376 173936
rect 137428 173924 137434 173936
rect 186314 173924 186320 173936
rect 137428 173896 186320 173924
rect 137428 173884 137434 173896
rect 186314 173884 186320 173896
rect 186372 173884 186378 173936
rect 411254 173884 411260 173936
rect 411312 173924 411318 173936
rect 424318 173924 424324 173936
rect 411312 173896 424324 173924
rect 411312 173884 411318 173896
rect 424318 173884 424324 173896
rect 424376 173884 424382 173936
rect 138750 172524 138756 172576
rect 138808 172564 138814 172576
rect 186314 172564 186320 172576
rect 138808 172536 186320 172564
rect 138808 172524 138814 172536
rect 186314 172524 186320 172536
rect 186372 172524 186378 172576
rect 411254 172524 411260 172576
rect 411312 172564 411318 172576
rect 421742 172564 421748 172576
rect 411312 172536 421748 172564
rect 411312 172524 411318 172536
rect 421742 172524 421748 172536
rect 421800 172524 421806 172576
rect 145834 171096 145840 171148
rect 145892 171136 145898 171148
rect 186314 171136 186320 171148
rect 145892 171108 186320 171136
rect 145892 171096 145898 171108
rect 186314 171096 186320 171108
rect 186372 171096 186378 171148
rect 166258 169736 166264 169788
rect 166316 169776 166322 169788
rect 186314 169776 186320 169788
rect 166316 169748 186320 169776
rect 166316 169736 166322 169748
rect 186314 169736 186320 169748
rect 186372 169736 186378 169788
rect 411254 169736 411260 169788
rect 411312 169776 411318 169788
rect 418982 169776 418988 169788
rect 411312 169748 418988 169776
rect 411312 169736 411318 169748
rect 418982 169736 418988 169748
rect 419040 169736 419046 169788
rect 136174 168376 136180 168428
rect 136232 168416 136238 168428
rect 186314 168416 186320 168428
rect 136232 168388 186320 168416
rect 136232 168376 136238 168388
rect 186314 168376 186320 168388
rect 186372 168376 186378 168428
rect 411254 168376 411260 168428
rect 411312 168416 411318 168428
rect 420270 168416 420276 168428
rect 411312 168388 420276 168416
rect 411312 168376 411318 168388
rect 420270 168376 420276 168388
rect 420328 168376 420334 168428
rect 138842 167084 138848 167136
rect 138900 167124 138906 167136
rect 186314 167124 186320 167136
rect 138900 167096 186320 167124
rect 138900 167084 138906 167096
rect 186314 167084 186320 167096
rect 186372 167084 186378 167136
rect 131942 167016 131948 167068
rect 132000 167056 132006 167068
rect 186406 167056 186412 167068
rect 132000 167028 186412 167056
rect 132000 167016 132006 167028
rect 186406 167016 186412 167028
rect 186464 167016 186470 167068
rect 164878 165588 164884 165640
rect 164936 165628 164942 165640
rect 186314 165628 186320 165640
rect 164936 165600 186320 165628
rect 164936 165588 164942 165600
rect 186314 165588 186320 165600
rect 186372 165588 186378 165640
rect 411254 165588 411260 165640
rect 411312 165628 411318 165640
rect 417418 165628 417424 165640
rect 411312 165600 417424 165628
rect 411312 165588 411318 165600
rect 417418 165588 417424 165600
rect 417476 165588 417482 165640
rect 138934 164228 138940 164280
rect 138992 164268 138998 164280
rect 186314 164268 186320 164280
rect 138992 164240 186320 164268
rect 138992 164228 138998 164240
rect 186314 164228 186320 164240
rect 186372 164228 186378 164280
rect 411254 164228 411260 164280
rect 411312 164268 411318 164280
rect 420178 164268 420184 164280
rect 411312 164240 420184 164268
rect 411312 164228 411318 164240
rect 420178 164228 420184 164240
rect 420236 164228 420242 164280
rect 132034 162868 132040 162920
rect 132092 162908 132098 162920
rect 186314 162908 186320 162920
rect 132092 162880 186320 162908
rect 132092 162868 132098 162880
rect 186314 162868 186320 162880
rect 186372 162868 186378 162920
rect 162118 161508 162124 161560
rect 162176 161548 162182 161560
rect 186314 161548 186320 161560
rect 162176 161520 186320 161548
rect 162176 161508 162182 161520
rect 186314 161508 186320 161520
rect 186372 161508 186378 161560
rect 135070 161440 135076 161492
rect 135128 161480 135134 161492
rect 186406 161480 186412 161492
rect 135128 161452 186412 161480
rect 135128 161440 135134 161452
rect 186406 161440 186412 161452
rect 186464 161440 186470 161492
rect 411254 161440 411260 161492
rect 411312 161480 411318 161492
rect 417602 161480 417608 161492
rect 411312 161452 417608 161480
rect 411312 161440 411318 161452
rect 417602 161440 417608 161452
rect 417660 161440 417666 161492
rect 136266 160080 136272 160132
rect 136324 160120 136330 160132
rect 186314 160120 186320 160132
rect 136324 160092 186320 160120
rect 136324 160080 136330 160092
rect 186314 160080 186320 160092
rect 186372 160080 186378 160132
rect 411254 160080 411260 160132
rect 411312 160120 411318 160132
rect 420362 160120 420368 160132
rect 411312 160092 420368 160120
rect 411312 160080 411318 160092
rect 420362 160080 420368 160092
rect 420420 160080 420426 160132
rect 132126 158720 132132 158772
rect 132184 158760 132190 158772
rect 186314 158760 186320 158772
rect 132184 158732 186320 158760
rect 132184 158720 132190 158732
rect 186314 158720 186320 158732
rect 186372 158720 186378 158772
rect 411254 158720 411260 158772
rect 411312 158760 411318 158772
rect 417510 158760 417516 158772
rect 411312 158732 417516 158760
rect 411312 158720 411318 158732
rect 417510 158720 417516 158732
rect 417568 158720 417574 158772
rect 139026 157360 139032 157412
rect 139084 157400 139090 157412
rect 186314 157400 186320 157412
rect 139084 157372 186320 157400
rect 139084 157360 139090 157372
rect 186314 157360 186320 157372
rect 186372 157360 186378 157412
rect 160738 155932 160744 155984
rect 160796 155972 160802 155984
rect 186314 155972 186320 155984
rect 160796 155944 186320 155972
rect 160796 155932 160802 155944
rect 186314 155932 186320 155944
rect 186372 155932 186378 155984
rect 411254 155932 411260 155984
rect 411312 155972 411318 155984
rect 419074 155972 419080 155984
rect 411312 155944 419080 155972
rect 411312 155932 411318 155944
rect 419074 155932 419080 155944
rect 419132 155932 419138 155984
rect 137462 154640 137468 154692
rect 137520 154680 137526 154692
rect 186314 154680 186320 154692
rect 137520 154652 186320 154680
rect 137520 154640 137526 154652
rect 186314 154640 186320 154652
rect 186372 154640 186378 154692
rect 133782 154572 133788 154624
rect 133840 154612 133846 154624
rect 186406 154612 186412 154624
rect 133840 154584 186412 154612
rect 133840 154572 133846 154584
rect 186406 154572 186412 154584
rect 186464 154572 186470 154624
rect 411254 154572 411260 154624
rect 411312 154612 411318 154624
rect 417694 154612 417700 154624
rect 411312 154584 417700 154612
rect 411312 154572 411318 154584
rect 417694 154572 417700 154584
rect 417752 154572 417758 154624
rect 145926 153212 145932 153264
rect 145984 153252 145990 153264
rect 186314 153252 186320 153264
rect 145984 153224 186320 153252
rect 145984 153212 145990 153224
rect 186314 153212 186320 153224
rect 186372 153212 186378 153264
rect 147122 151784 147128 151836
rect 147180 151824 147186 151836
rect 186314 151824 186320 151836
rect 147180 151796 186320 151824
rect 147180 151784 147186 151796
rect 186314 151784 186320 151796
rect 186372 151784 186378 151836
rect 411254 151784 411260 151836
rect 411312 151824 411318 151836
rect 414934 151824 414940 151836
rect 411312 151796 414940 151824
rect 411312 151784 411318 151796
rect 414934 151784 414940 151796
rect 414992 151784 414998 151836
rect 146018 150424 146024 150476
rect 146076 150464 146082 150476
rect 186314 150464 186320 150476
rect 146076 150436 186320 150464
rect 146076 150424 146082 150436
rect 186314 150424 186320 150436
rect 186372 150424 186378 150476
rect 411254 150424 411260 150476
rect 411312 150464 411318 150476
rect 417786 150464 417792 150476
rect 411312 150436 417792 150464
rect 411312 150424 411318 150436
rect 417786 150424 417792 150436
rect 417844 150424 417850 150476
rect 144178 149132 144184 149184
rect 144236 149172 144242 149184
rect 186314 149172 186320 149184
rect 144236 149144 186320 149172
rect 144236 149132 144242 149144
rect 186314 149132 186320 149144
rect 186372 149132 186378 149184
rect 137554 149064 137560 149116
rect 137612 149104 137618 149116
rect 186406 149104 186412 149116
rect 137612 149076 186412 149104
rect 137612 149064 137618 149076
rect 186406 149064 186412 149076
rect 186464 149064 186470 149116
rect 132218 147636 132224 147688
rect 132276 147676 132282 147688
rect 186314 147676 186320 147688
rect 132276 147648 186320 147676
rect 132276 147636 132282 147648
rect 186314 147636 186320 147648
rect 186372 147636 186378 147688
rect 411254 147636 411260 147688
rect 411312 147676 411318 147688
rect 415026 147676 415032 147688
rect 411312 147648 415032 147676
rect 411312 147636 411318 147648
rect 415026 147636 415032 147648
rect 415084 147636 415090 147688
rect 144270 146276 144276 146328
rect 144328 146316 144334 146328
rect 186314 146316 186320 146328
rect 144328 146288 186320 146316
rect 144328 146276 144334 146288
rect 186314 146276 186320 146288
rect 186372 146276 186378 146328
rect 411254 146276 411260 146328
rect 411312 146316 411318 146328
rect 421834 146316 421840 146328
rect 411312 146288 421840 146316
rect 411312 146276 411318 146288
rect 421834 146276 421840 146288
rect 421892 146276 421898 146328
rect 143074 144916 143080 144968
rect 143132 144956 143138 144968
rect 186314 144956 186320 144968
rect 143132 144928 186320 144956
rect 143132 144916 143138 144928
rect 186314 144916 186320 144928
rect 186372 144916 186378 144968
rect 411254 144916 411260 144968
rect 411312 144956 411318 144968
rect 417878 144956 417884 144968
rect 411312 144928 417884 144956
rect 411312 144916 411318 144928
rect 417878 144916 417884 144928
rect 417936 144916 417942 144968
rect 141602 143556 141608 143608
rect 141660 143596 141666 143608
rect 186314 143596 186320 143608
rect 141660 143568 186320 143596
rect 141660 143556 141666 143568
rect 186314 143556 186320 143568
rect 186372 143556 186378 143608
rect 144362 142196 144368 142248
rect 144420 142236 144426 142248
rect 186406 142236 186412 142248
rect 144420 142208 186412 142236
rect 144420 142196 144426 142208
rect 186406 142196 186412 142208
rect 186464 142196 186470 142248
rect 142982 142128 142988 142180
rect 143040 142168 143046 142180
rect 186314 142168 186320 142180
rect 143040 142140 186320 142168
rect 143040 142128 143046 142140
rect 186314 142128 186320 142140
rect 186372 142128 186378 142180
rect 411254 142128 411260 142180
rect 411312 142168 411318 142180
rect 429930 142168 429936 142180
rect 411312 142140 429936 142168
rect 411312 142128 411318 142140
rect 429930 142128 429936 142140
rect 429988 142128 429994 142180
rect 411254 140768 411260 140820
rect 411312 140808 411318 140820
rect 421926 140808 421932 140820
rect 411312 140780 421932 140808
rect 411312 140768 411318 140780
rect 421926 140768 421932 140780
rect 421984 140768 421990 140820
rect 137646 139408 137652 139460
rect 137704 139448 137710 139460
rect 186314 139448 186320 139460
rect 137704 139420 186320 139448
rect 137704 139408 137710 139420
rect 186314 139408 186320 139420
rect 186372 139408 186378 139460
rect 414658 139340 414664 139392
rect 414716 139380 414722 139392
rect 580166 139380 580172 139392
rect 414716 139352 580172 139380
rect 414716 139340 414722 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 143166 137980 143172 138032
rect 143224 138020 143230 138032
rect 186314 138020 186320 138032
rect 143224 137992 186320 138020
rect 143224 137980 143230 137992
rect 186314 137980 186320 137992
rect 186372 137980 186378 138032
rect 411254 137980 411260 138032
rect 411312 138020 411318 138032
rect 431310 138020 431316 138032
rect 411312 137992 431316 138020
rect 411312 137980 411318 137992
rect 431310 137980 431316 137992
rect 431368 137980 431374 138032
rect 141694 136620 141700 136672
rect 141752 136660 141758 136672
rect 186314 136660 186320 136672
rect 141752 136632 186320 136660
rect 141752 136620 141758 136632
rect 186314 136620 186320 136632
rect 186372 136620 186378 136672
rect 411254 136620 411260 136672
rect 411312 136660 411318 136672
rect 422018 136660 422024 136672
rect 411312 136632 422024 136660
rect 411312 136620 411318 136632
rect 422018 136620 422024 136632
rect 422076 136620 422082 136672
rect 143258 135328 143264 135380
rect 143316 135368 143322 135380
rect 186314 135368 186320 135380
rect 143316 135340 186320 135368
rect 143316 135328 143322 135340
rect 186314 135328 186320 135340
rect 186372 135328 186378 135380
rect 137738 135260 137744 135312
rect 137796 135300 137802 135312
rect 186406 135300 186412 135312
rect 137796 135272 186412 135300
rect 137796 135260 137802 135272
rect 186406 135260 186412 135272
rect 186464 135260 186470 135312
rect 140406 133900 140412 133952
rect 140464 133940 140470 133952
rect 186314 133940 186320 133952
rect 140464 133912 186320 133940
rect 140464 133900 140470 133912
rect 186314 133900 186320 133912
rect 186372 133900 186378 133952
rect 411254 133900 411260 133952
rect 411312 133940 411318 133952
rect 432690 133940 432696 133952
rect 411312 133912 432696 133940
rect 411312 133900 411318 133912
rect 432690 133900 432696 133912
rect 432748 133900 432754 133952
rect 137830 132472 137836 132524
rect 137888 132512 137894 132524
rect 186314 132512 186320 132524
rect 137888 132484 186320 132512
rect 137888 132472 137894 132484
rect 186314 132472 186320 132484
rect 186372 132472 186378 132524
rect 411254 132472 411260 132524
rect 411312 132512 411318 132524
rect 420454 132512 420460 132524
rect 411312 132484 420460 132512
rect 411312 132472 411318 132484
rect 420454 132472 420460 132484
rect 420512 132472 420518 132524
rect 103330 132268 103336 132320
rect 103388 132308 103394 132320
rect 133138 132308 133144 132320
rect 103388 132280 133144 132308
rect 103388 132268 103394 132280
rect 133138 132268 133144 132280
rect 133196 132268 133202 132320
rect 100662 132200 100668 132252
rect 100720 132240 100726 132252
rect 131666 132240 131672 132252
rect 100720 132212 131672 132240
rect 100720 132200 100726 132212
rect 131666 132200 131672 132212
rect 131724 132200 131730 132252
rect 97718 132132 97724 132184
rect 97776 132172 97782 132184
rect 130562 132172 130568 132184
rect 97776 132144 130568 132172
rect 97776 132132 97782 132144
rect 130562 132132 130568 132144
rect 130620 132132 130626 132184
rect 108942 132064 108948 132116
rect 109000 132104 109006 132116
rect 188706 132104 188712 132116
rect 109000 132076 188712 132104
rect 109000 132064 109006 132076
rect 188706 132064 188712 132076
rect 188764 132064 188770 132116
rect 97810 131996 97816 132048
rect 97868 132036 97874 132048
rect 188982 132036 188988 132048
rect 97868 132008 188988 132036
rect 97868 131996 97874 132008
rect 188982 131996 188988 132008
rect 189040 131996 189046 132048
rect 88242 131928 88248 131980
rect 88300 131968 88306 131980
rect 182818 131968 182824 131980
rect 88300 131940 182824 131968
rect 88300 131928 88306 131940
rect 182818 131928 182824 131940
rect 182876 131928 182882 131980
rect 92382 131860 92388 131912
rect 92440 131900 92446 131912
rect 188798 131900 188804 131912
rect 92440 131872 188804 131900
rect 92440 131860 92446 131872
rect 188798 131860 188804 131872
rect 188856 131860 188862 131912
rect 92290 131792 92296 131844
rect 92348 131832 92354 131844
rect 188890 131832 188896 131844
rect 92348 131804 188896 131832
rect 92348 131792 92354 131804
rect 188890 131792 188896 131804
rect 188948 131792 188954 131844
rect 48222 131724 48228 131776
rect 48280 131764 48286 131776
rect 188614 131764 188620 131776
rect 48280 131736 188620 131764
rect 48280 131724 48286 131736
rect 188614 131724 188620 131736
rect 188672 131724 188678 131776
rect 419350 131452 419356 131504
rect 419408 131492 419414 131504
rect 534626 131492 534632 131504
rect 419408 131464 534632 131492
rect 419408 131452 419414 131464
rect 534626 131452 534632 131464
rect 534684 131452 534690 131504
rect 410518 131384 410524 131436
rect 410576 131424 410582 131436
rect 444650 131424 444656 131436
rect 410576 131396 444656 131424
rect 410576 131384 410582 131396
rect 444650 131384 444656 131396
rect 444708 131384 444714 131436
rect 414658 131316 414664 131368
rect 414716 131356 414722 131368
rect 484578 131356 484584 131368
rect 414716 131328 484584 131356
rect 414716 131316 414722 131328
rect 484578 131316 484584 131328
rect 484636 131316 484642 131368
rect 414750 131248 414756 131300
rect 414808 131288 414814 131300
rect 494606 131288 494612 131300
rect 414808 131260 494612 131288
rect 414808 131248 414814 131260
rect 494606 131248 494612 131260
rect 494664 131248 494670 131300
rect 1302 131180 1308 131232
rect 1360 131220 1366 131232
rect 55122 131220 55128 131232
rect 1360 131192 55128 131220
rect 1360 131180 1366 131192
rect 55122 131180 55128 131192
rect 55180 131180 55186 131232
rect 414842 131180 414848 131232
rect 414900 131220 414906 131232
rect 504634 131220 504640 131232
rect 414900 131192 504640 131220
rect 414900 131180 414906 131192
rect 504634 131180 504640 131192
rect 504692 131180 504698 131232
rect 2682 131112 2688 131164
rect 2740 131152 2746 131164
rect 104894 131152 104900 131164
rect 2740 131124 104900 131152
rect 2740 131112 2746 131124
rect 104894 131112 104900 131124
rect 104952 131112 104958 131164
rect 141878 131112 141884 131164
rect 141936 131152 141942 131164
rect 186314 131152 186320 131164
rect 141936 131124 186320 131152
rect 141936 131112 141942 131124
rect 186314 131112 186320 131124
rect 186372 131112 186378 131164
rect 96522 130704 96528 130756
rect 96580 130744 96586 130756
rect 130654 130744 130660 130756
rect 96580 130716 130660 130744
rect 96580 130704 96586 130716
rect 130654 130704 130660 130716
rect 130712 130704 130718 130756
rect 85482 130636 85488 130688
rect 85540 130676 85546 130688
rect 188246 130676 188252 130688
rect 85540 130648 188252 130676
rect 85540 130636 85546 130648
rect 188246 130636 188252 130648
rect 188304 130636 188310 130688
rect 85390 130568 85396 130620
rect 85448 130608 85454 130620
rect 188154 130608 188160 130620
rect 85448 130580 188160 130608
rect 85448 130568 85454 130580
rect 188154 130568 188160 130580
rect 188212 130568 188218 130620
rect 86862 130500 86868 130552
rect 86920 130540 86926 130552
rect 189810 130540 189816 130552
rect 86920 130512 189816 130540
rect 86920 130500 86926 130512
rect 189810 130500 189816 130512
rect 189868 130500 189874 130552
rect 85298 130432 85304 130484
rect 85356 130472 85362 130484
rect 189718 130472 189724 130484
rect 85356 130444 189724 130472
rect 85356 130432 85362 130444
rect 189718 130432 189724 130444
rect 189776 130432 189782 130484
rect 84102 130364 84108 130416
rect 84160 130404 84166 130416
rect 189810 130404 189816 130416
rect 84160 130376 189816 130404
rect 84160 130364 84166 130376
rect 189810 130364 189816 130376
rect 189868 130364 189874 130416
rect 434622 130364 434628 130416
rect 434680 130404 434686 130416
rect 454586 130404 454592 130416
rect 434680 130376 454592 130404
rect 434680 130364 434686 130376
rect 454586 130364 454592 130376
rect 454644 130364 454650 130416
rect 418890 130024 418896 130076
rect 418948 130064 418954 130076
rect 474734 130064 474740 130076
rect 418948 130036 474740 130064
rect 418948 130024 418954 130036
rect 474734 130024 474740 130036
rect 474792 130024 474798 130076
rect 413278 129956 413284 130008
rect 413336 129996 413342 130008
rect 514754 129996 514760 130008
rect 413336 129968 514760 129996
rect 413336 129956 413342 129968
rect 514754 129956 514760 129968
rect 514812 129956 514818 130008
rect 413462 129888 413468 129940
rect 413520 129928 413526 129940
rect 524598 129928 524604 129940
rect 413520 129900 524604 129928
rect 413520 129888 413526 129900
rect 524598 129888 524604 129900
rect 524656 129888 524662 129940
rect 415210 129820 415216 129872
rect 415268 129860 415274 129872
rect 539318 129860 539324 129872
rect 415268 129832 539324 129860
rect 415268 129820 415274 129832
rect 539318 129820 539324 129832
rect 539376 129820 539382 129872
rect 144454 129752 144460 129804
rect 144512 129792 144518 129804
rect 186314 129792 186320 129804
rect 144512 129764 186320 129792
rect 144512 129752 144518 129764
rect 186314 129752 186320 129764
rect 186372 129752 186378 129804
rect 413370 129752 413376 129804
rect 413428 129792 413434 129804
rect 542446 129792 542452 129804
rect 413428 129764 542452 129792
rect 413428 129752 413434 129764
rect 542446 129752 542452 129764
rect 542504 129752 542510 129804
rect 131114 129684 131120 129736
rect 131172 129724 131178 129736
rect 169018 129724 169024 129736
rect 131172 129696 169024 129724
rect 131172 129684 131178 129696
rect 169018 129684 169024 129696
rect 169076 129684 169082 129736
rect 131206 129616 131212 129668
rect 131264 129656 131270 129668
rect 159358 129656 159364 129668
rect 131264 129628 159364 129656
rect 131264 129616 131270 129628
rect 159358 129616 159364 129628
rect 159416 129616 159422 129668
rect 411254 128460 411260 128512
rect 411312 128500 411318 128512
rect 420546 128500 420552 128512
rect 411312 128472 420552 128500
rect 411312 128460 411318 128472
rect 420546 128460 420552 128472
rect 420604 128460 420610 128512
rect 425790 128460 425796 128512
rect 425848 128500 425854 128512
rect 434622 128500 434628 128512
rect 425848 128472 434628 128500
rect 425848 128460 425854 128472
rect 434622 128460 434628 128472
rect 434680 128460 434686 128512
rect 419258 128392 419264 128444
rect 419316 128432 419322 128444
rect 437474 128432 437480 128444
rect 419316 128404 437480 128432
rect 419316 128392 419322 128404
rect 437474 128392 437480 128404
rect 437532 128392 437538 128444
rect 141786 128324 141792 128376
rect 141844 128364 141850 128376
rect 186314 128364 186320 128376
rect 141844 128336 186320 128364
rect 141844 128324 141850 128336
rect 186314 128324 186320 128336
rect 186372 128324 186378 128376
rect 412450 128324 412456 128376
rect 412508 128364 412514 128376
rect 542354 128364 542360 128376
rect 412508 128336 542360 128364
rect 412508 128324 412514 128336
rect 542354 128324 542360 128336
rect 542412 128324 542418 128376
rect 131206 128256 131212 128308
rect 131264 128296 131270 128308
rect 142798 128296 142804 128308
rect 131264 128268 142804 128296
rect 131264 128256 131270 128268
rect 142798 128256 142804 128268
rect 142856 128256 142862 128308
rect 131758 128188 131764 128240
rect 131816 128228 131822 128240
rect 135990 128228 135996 128240
rect 131816 128200 135996 128228
rect 131816 128188 131822 128200
rect 135990 128188 135996 128200
rect 136048 128188 136054 128240
rect 411254 127032 411260 127084
rect 411312 127072 411318 127084
rect 435450 127072 435456 127084
rect 411312 127044 435456 127072
rect 411312 127032 411318 127044
rect 435450 127032 435456 127044
rect 435508 127032 435514 127084
rect 140498 126964 140504 127016
rect 140556 127004 140562 127016
rect 186314 127004 186320 127016
rect 140556 126976 186320 127004
rect 140556 126964 140562 126976
rect 186314 126964 186320 126976
rect 186372 126964 186378 127016
rect 413830 126964 413836 127016
rect 413888 127004 413894 127016
rect 437474 127004 437480 127016
rect 413888 126976 437480 127004
rect 413888 126964 413894 126976
rect 437474 126964 437480 126976
rect 437532 126964 437538 127016
rect 131114 126896 131120 126948
rect 131172 126936 131178 126948
rect 157978 126936 157984 126948
rect 131172 126908 157984 126936
rect 131172 126896 131178 126908
rect 157978 126896 157984 126908
rect 158036 126896 158042 126948
rect 131206 126828 131212 126880
rect 131264 126868 131270 126880
rect 135898 126868 135904 126880
rect 131264 126840 135904 126868
rect 131264 126828 131270 126840
rect 135898 126828 135904 126840
rect 135956 126828 135962 126880
rect 131114 125672 131120 125724
rect 131172 125712 131178 125724
rect 134518 125712 134524 125724
rect 131172 125684 134524 125712
rect 131172 125672 131178 125684
rect 134518 125672 134524 125684
rect 134576 125672 134582 125724
rect 144546 125604 144552 125656
rect 144604 125644 144610 125656
rect 186314 125644 186320 125656
rect 144604 125616 186320 125644
rect 144604 125604 144610 125616
rect 186314 125604 186320 125616
rect 186372 125604 186378 125656
rect 413738 125604 413744 125656
rect 413796 125644 413802 125656
rect 437474 125644 437480 125656
rect 413796 125616 437480 125644
rect 413796 125604 413802 125616
rect 437474 125604 437480 125616
rect 437532 125604 437538 125656
rect 131206 125536 131212 125588
rect 131264 125576 131270 125588
rect 186958 125576 186964 125588
rect 131264 125548 186964 125576
rect 131264 125536 131270 125548
rect 186958 125536 186964 125548
rect 187016 125536 187022 125588
rect 131574 125468 131580 125520
rect 131632 125508 131638 125520
rect 141418 125508 141424 125520
rect 131632 125480 141424 125508
rect 131632 125468 131638 125480
rect 141418 125468 141424 125480
rect 141476 125468 141482 125520
rect 411254 124244 411260 124296
rect 411312 124284 411318 124296
rect 416222 124284 416228 124296
rect 411312 124256 416228 124284
rect 411312 124244 411318 124256
rect 416222 124244 416228 124256
rect 416280 124244 416286 124296
rect 141970 124176 141976 124228
rect 142028 124216 142034 124228
rect 186314 124216 186320 124228
rect 142028 124188 186320 124216
rect 142028 124176 142034 124188
rect 186314 124176 186320 124188
rect 186372 124176 186378 124228
rect 413646 124176 413652 124228
rect 413704 124216 413710 124228
rect 437474 124216 437480 124228
rect 413704 124188 437480 124216
rect 413704 124176 413710 124188
rect 437474 124176 437480 124188
rect 437532 124176 437538 124228
rect 131758 124108 131764 124160
rect 131816 124148 131822 124160
rect 156598 124148 156604 124160
rect 131816 124120 156604 124148
rect 131816 124108 131822 124120
rect 156598 124108 156604 124120
rect 156656 124108 156662 124160
rect 131114 124040 131120 124092
rect 131172 124080 131178 124092
rect 136082 124080 136088 124092
rect 131172 124052 136088 124080
rect 131172 124040 131178 124052
rect 136082 124040 136088 124052
rect 136140 124040 136146 124092
rect 411254 122884 411260 122936
rect 411312 122924 411318 122936
rect 428550 122924 428556 122936
rect 411312 122896 428556 122924
rect 411312 122884 411318 122896
rect 428550 122884 428556 122896
rect 428608 122884 428614 122936
rect 144638 122816 144644 122868
rect 144696 122856 144702 122868
rect 186314 122856 186320 122868
rect 144696 122828 186320 122856
rect 144696 122816 144702 122828
rect 186314 122816 186320 122828
rect 186372 122816 186378 122868
rect 413554 122816 413560 122868
rect 413612 122856 413618 122868
rect 437474 122856 437480 122868
rect 413612 122828 437480 122856
rect 413612 122816 413618 122828
rect 437474 122816 437480 122828
rect 437532 122816 437538 122868
rect 131114 122748 131120 122800
rect 131172 122788 131178 122800
rect 155218 122788 155224 122800
rect 131172 122760 155224 122788
rect 131172 122748 131178 122760
rect 155218 122748 155224 122760
rect 155276 122748 155282 122800
rect 131206 122680 131212 122732
rect 131264 122720 131270 122732
rect 141510 122720 141516 122732
rect 131264 122692 141516 122720
rect 131264 122680 131270 122692
rect 141510 122680 141516 122692
rect 141568 122680 141574 122732
rect 131482 122612 131488 122664
rect 131540 122652 131546 122664
rect 133230 122652 133236 122664
rect 131540 122624 133236 122652
rect 131540 122612 131546 122624
rect 133230 122612 133236 122624
rect 133288 122612 133294 122664
rect 423766 121524 423772 121576
rect 423824 121564 423830 121576
rect 425790 121564 425796 121576
rect 423824 121536 425796 121564
rect 423824 121524 423830 121536
rect 425790 121524 425796 121536
rect 425848 121524 425854 121576
rect 141418 121456 141424 121508
rect 141476 121496 141482 121508
rect 186314 121496 186320 121508
rect 141476 121468 186320 121496
rect 141476 121456 141482 121468
rect 186314 121456 186320 121468
rect 186372 121456 186378 121508
rect 131206 121388 131212 121440
rect 131264 121428 131270 121440
rect 187050 121428 187056 121440
rect 131264 121400 187056 121428
rect 131264 121388 131270 121400
rect 187050 121388 187056 121400
rect 187108 121388 187114 121440
rect 131114 121320 131120 121372
rect 131172 121360 131178 121372
rect 142890 121360 142896 121372
rect 131172 121332 142896 121360
rect 131172 121320 131178 121332
rect 142890 121320 142896 121332
rect 142948 121320 142954 121372
rect 410610 120708 410616 120760
rect 410668 120748 410674 120760
rect 423766 120748 423772 120760
rect 410668 120720 423772 120748
rect 410668 120708 410674 120720
rect 423766 120708 423772 120720
rect 423824 120708 423830 120760
rect 411254 120096 411260 120148
rect 411312 120136 411318 120148
rect 436830 120136 436836 120148
rect 411312 120108 436836 120136
rect 411312 120096 411318 120108
rect 436830 120096 436836 120108
rect 436888 120096 436894 120148
rect 131114 120028 131120 120080
rect 131172 120068 131178 120080
rect 152458 120068 152464 120080
rect 131172 120040 152464 120068
rect 131172 120028 131178 120040
rect 152458 120028 152464 120040
rect 152516 120028 152522 120080
rect 132310 119960 132316 120012
rect 132368 120000 132374 120012
rect 134610 120000 134616 120012
rect 132368 119972 134616 120000
rect 132368 119960 132374 119972
rect 134610 119960 134616 119972
rect 134668 119960 134674 120012
rect 142798 118668 142804 118720
rect 142856 118708 142862 118720
rect 186314 118708 186320 118720
rect 142856 118680 186320 118708
rect 142856 118668 142862 118680
rect 186314 118668 186320 118680
rect 186372 118668 186378 118720
rect 411254 118668 411260 118720
rect 411312 118708 411318 118720
rect 416314 118708 416320 118720
rect 411312 118680 416320 118708
rect 411312 118668 411318 118680
rect 416314 118668 416320 118680
rect 416372 118668 416378 118720
rect 131298 118600 131304 118652
rect 131356 118640 131362 118652
rect 151078 118640 151084 118652
rect 131356 118612 151084 118640
rect 131356 118600 131362 118612
rect 151078 118600 151084 118612
rect 151136 118600 151142 118652
rect 131206 118532 131212 118584
rect 131264 118572 131270 118584
rect 134702 118572 134708 118584
rect 131264 118544 134708 118572
rect 131264 118532 131270 118544
rect 134702 118532 134708 118544
rect 134760 118532 134766 118584
rect 131114 118464 131120 118516
rect 131172 118504 131178 118516
rect 134794 118504 134800 118516
rect 131172 118476 134800 118504
rect 131172 118464 131178 118476
rect 134794 118464 134800 118476
rect 134852 118464 134858 118516
rect 134610 117376 134616 117428
rect 134668 117416 134674 117428
rect 186406 117416 186412 117428
rect 134668 117388 186412 117416
rect 134668 117376 134674 117388
rect 186406 117376 186412 117388
rect 186464 117376 186470 117428
rect 131850 117308 131856 117360
rect 131908 117348 131914 117360
rect 186314 117348 186320 117360
rect 131908 117320 186320 117348
rect 131908 117308 131914 117320
rect 186314 117308 186320 117320
rect 186372 117308 186378 117360
rect 131206 117240 131212 117292
rect 131264 117280 131270 117292
rect 148318 117280 148324 117292
rect 131264 117252 148324 117280
rect 131264 117240 131270 117252
rect 148318 117240 148324 117252
rect 148376 117240 148382 117292
rect 131114 117172 131120 117224
rect 131172 117212 131178 117224
rect 134886 117212 134892 117224
rect 131172 117184 134892 117212
rect 131172 117172 131178 117184
rect 134886 117172 134892 117184
rect 134944 117172 134950 117224
rect 142890 115948 142896 116000
rect 142948 115988 142954 116000
rect 186314 115988 186320 116000
rect 142948 115960 186320 115988
rect 142948 115948 142954 115960
rect 186314 115948 186320 115960
rect 186372 115948 186378 116000
rect 132310 115880 132316 115932
rect 132368 115920 132374 115932
rect 145558 115920 145564 115932
rect 132368 115892 145564 115920
rect 132368 115880 132374 115892
rect 145558 115880 145564 115892
rect 145616 115880 145622 115932
rect 131206 115472 131212 115524
rect 131264 115512 131270 115524
rect 134978 115512 134984 115524
rect 131264 115484 134984 115512
rect 131264 115472 131270 115484
rect 134978 115472 134984 115484
rect 135036 115472 135042 115524
rect 134518 114520 134524 114572
rect 134576 114560 134582 114572
rect 186314 114560 186320 114572
rect 134576 114532 186320 114560
rect 134576 114520 134582 114532
rect 186314 114520 186320 114532
rect 186372 114520 186378 114572
rect 411254 114520 411260 114572
rect 411312 114560 411318 114572
rect 419166 114560 419172 114572
rect 411312 114532 419172 114560
rect 411312 114520 411318 114532
rect 419166 114520 419172 114532
rect 419224 114520 419230 114572
rect 131298 114452 131304 114504
rect 131356 114492 131362 114504
rect 147030 114492 147036 114504
rect 131356 114464 147036 114492
rect 131356 114452 131362 114464
rect 147030 114452 147036 114464
rect 147088 114452 147094 114504
rect 411898 114452 411904 114504
rect 411956 114492 411962 114504
rect 437474 114492 437480 114504
rect 411956 114464 437480 114492
rect 411956 114452 411962 114464
rect 437474 114452 437480 114464
rect 437532 114452 437538 114504
rect 131206 114384 131212 114436
rect 131264 114424 131270 114436
rect 146938 114424 146944 114436
rect 131264 114396 146944 114424
rect 131264 114384 131270 114396
rect 146938 114384 146944 114396
rect 146996 114384 147002 114436
rect 131114 114316 131120 114368
rect 131172 114356 131178 114368
rect 133322 114356 133328 114368
rect 131172 114328 133328 114356
rect 131172 114316 131178 114328
rect 133322 114316 133328 114328
rect 133380 114316 133386 114368
rect 131666 113160 131672 113212
rect 131724 113200 131730 113212
rect 186314 113200 186320 113212
rect 131724 113172 186320 113200
rect 131724 113160 131730 113172
rect 186314 113160 186320 113172
rect 186372 113160 186378 113212
rect 411254 113160 411260 113212
rect 411312 113200 411318 113212
rect 416406 113200 416412 113212
rect 411312 113172 416412 113200
rect 411312 113160 411318 113172
rect 416406 113160 416412 113172
rect 416464 113160 416470 113212
rect 131206 113092 131212 113144
rect 131264 113132 131270 113144
rect 145650 113132 145656 113144
rect 131264 113104 145656 113132
rect 131264 113092 131270 113104
rect 145650 113092 145656 113104
rect 145708 113092 145714 113144
rect 412082 113092 412088 113144
rect 412140 113132 412146 113144
rect 437474 113132 437480 113144
rect 412140 113104 437480 113132
rect 412140 113092 412146 113104
rect 437474 113092 437480 113104
rect 437532 113092 437538 113144
rect 131114 113024 131120 113076
rect 131172 113064 131178 113076
rect 140130 113064 140136 113076
rect 131172 113036 140136 113064
rect 131172 113024 131178 113036
rect 140130 113024 140136 113036
rect 140188 113024 140194 113076
rect 135898 111868 135904 111920
rect 135956 111908 135962 111920
rect 186406 111908 186412 111920
rect 135956 111880 186412 111908
rect 135956 111868 135962 111880
rect 186406 111868 186412 111880
rect 186464 111868 186470 111920
rect 134702 111800 134708 111852
rect 134760 111840 134766 111852
rect 186314 111840 186320 111852
rect 134760 111812 186320 111840
rect 134760 111800 134766 111812
rect 186314 111800 186320 111812
rect 186372 111800 186378 111852
rect 131114 111732 131120 111784
rect 131172 111772 131178 111784
rect 140038 111772 140044 111784
rect 131172 111744 140044 111772
rect 131172 111732 131178 111744
rect 140038 111732 140044 111744
rect 140096 111732 140102 111784
rect 131206 111664 131212 111716
rect 131264 111704 131270 111716
rect 133414 111704 133420 111716
rect 131264 111676 133420 111704
rect 131264 111664 131270 111676
rect 133414 111664 133420 111676
rect 133472 111664 133478 111716
rect 131206 110372 131212 110424
rect 131264 110412 131270 110424
rect 187142 110412 187148 110424
rect 131264 110384 187148 110412
rect 131264 110372 131270 110384
rect 187142 110372 187148 110384
rect 187200 110372 187206 110424
rect 421558 110372 421564 110424
rect 421616 110412 421622 110424
rect 437474 110412 437480 110424
rect 421616 110384 437480 110412
rect 421616 110372 421622 110384
rect 437474 110372 437480 110384
rect 437532 110372 437538 110424
rect 131114 110304 131120 110356
rect 131172 110344 131178 110356
rect 145742 110344 145748 110356
rect 131172 110316 145748 110344
rect 131172 110304 131178 110316
rect 145742 110304 145748 110316
rect 145800 110304 145806 110356
rect 131206 110236 131212 110288
rect 131264 110276 131270 110288
rect 137278 110276 137284 110288
rect 131264 110248 137284 110276
rect 131264 110236 131270 110248
rect 137278 110236 137284 110248
rect 137336 110236 137342 110288
rect 135990 109012 135996 109064
rect 136048 109052 136054 109064
rect 186314 109052 186320 109064
rect 136048 109024 186320 109052
rect 136048 109012 136054 109024
rect 186314 109012 186320 109024
rect 186372 109012 186378 109064
rect 411254 109012 411260 109064
rect 411312 109052 411318 109064
rect 417970 109052 417976 109064
rect 411312 109024 417976 109052
rect 411312 109012 411318 109024
rect 417970 109012 417976 109024
rect 418028 109012 418034 109064
rect 131206 108944 131212 108996
rect 131264 108984 131270 108996
rect 140222 108984 140228 108996
rect 131264 108956 140228 108984
rect 131264 108944 131270 108956
rect 140222 108944 140228 108956
rect 140280 108944 140286 108996
rect 416038 108944 416044 108996
rect 416096 108984 416102 108996
rect 437474 108984 437480 108996
rect 416096 108956 437480 108984
rect 416096 108944 416102 108956
rect 437474 108944 437480 108956
rect 437532 108944 437538 108996
rect 131114 108876 131120 108928
rect 131172 108916 131178 108928
rect 133598 108916 133604 108928
rect 131172 108888 133604 108916
rect 131172 108876 131178 108888
rect 133598 108876 133604 108888
rect 133656 108876 133662 108928
rect 131666 108468 131672 108520
rect 131724 108508 131730 108520
rect 132310 108508 132316 108520
rect 131724 108480 132316 108508
rect 131724 108468 131730 108480
rect 132310 108468 132316 108480
rect 132368 108468 132374 108520
rect 131666 108332 131672 108384
rect 131724 108372 131730 108384
rect 132034 108372 132040 108384
rect 131724 108344 132040 108372
rect 131724 108332 131730 108344
rect 132034 108332 132040 108344
rect 132092 108332 132098 108384
rect 131574 108264 131580 108316
rect 131632 108304 131638 108316
rect 132126 108304 132132 108316
rect 131632 108276 132132 108304
rect 131632 108264 131638 108276
rect 132126 108264 132132 108276
rect 132184 108264 132190 108316
rect 133230 107652 133236 107704
rect 133288 107692 133294 107704
rect 186314 107692 186320 107704
rect 133288 107664 186320 107692
rect 133288 107652 133294 107664
rect 186314 107652 186320 107664
rect 186372 107652 186378 107704
rect 411254 107652 411260 107704
rect 411312 107692 411318 107704
rect 416498 107692 416504 107704
rect 411312 107664 416504 107692
rect 411312 107652 411318 107664
rect 416498 107652 416504 107664
rect 416556 107652 416562 107704
rect 131114 107584 131120 107636
rect 131172 107624 131178 107636
rect 133506 107624 133512 107636
rect 131172 107596 133512 107624
rect 131172 107584 131178 107596
rect 133506 107584 133512 107596
rect 133564 107584 133570 107636
rect 411990 107584 411996 107636
rect 412048 107624 412054 107636
rect 437474 107624 437480 107636
rect 412048 107596 437480 107624
rect 412048 107584 412054 107596
rect 437474 107584 437480 107596
rect 437532 107584 437538 107636
rect 131298 107516 131304 107568
rect 131356 107556 131362 107568
rect 138658 107556 138664 107568
rect 131356 107528 138664 107556
rect 131356 107516 131362 107528
rect 138658 107516 138664 107528
rect 138716 107516 138722 107568
rect 131206 107448 131212 107500
rect 131264 107488 131270 107500
rect 140314 107488 140320 107500
rect 131264 107460 140320 107488
rect 131264 107448 131270 107460
rect 140314 107448 140320 107460
rect 140372 107448 140378 107500
rect 140038 106292 140044 106344
rect 140096 106332 140102 106344
rect 186314 106332 186320 106344
rect 140096 106304 186320 106332
rect 140096 106292 140102 106304
rect 186314 106292 186320 106304
rect 186372 106292 186378 106344
rect 131114 106224 131120 106276
rect 131172 106264 131178 106276
rect 137370 106264 137376 106276
rect 131172 106236 137376 106264
rect 131172 106224 131178 106236
rect 137370 106224 137376 106236
rect 137428 106224 137434 106276
rect 131206 105952 131212 106004
rect 131264 105992 131270 106004
rect 133690 105992 133696 106004
rect 131264 105964 133696 105992
rect 131264 105952 131270 105964
rect 133690 105952 133696 105964
rect 133748 105952 133754 106004
rect 136082 104932 136088 104984
rect 136140 104972 136146 104984
rect 186406 104972 186412 104984
rect 136140 104944 186412 104972
rect 136140 104932 136146 104944
rect 186406 104932 186412 104944
rect 186464 104932 186470 104984
rect 134794 104864 134800 104916
rect 134852 104904 134858 104916
rect 186314 104904 186320 104916
rect 134852 104876 186320 104904
rect 134852 104864 134858 104876
rect 186314 104864 186320 104876
rect 186372 104864 186378 104916
rect 131206 104796 131212 104848
rect 131264 104836 131270 104848
rect 187234 104836 187240 104848
rect 131264 104808 187240 104836
rect 131264 104796 131270 104808
rect 187234 104796 187240 104808
rect 187292 104796 187298 104848
rect 421650 104796 421656 104848
rect 421708 104836 421714 104848
rect 437474 104836 437480 104848
rect 421708 104808 437480 104836
rect 421708 104796 421714 104808
rect 437474 104796 437480 104808
rect 437532 104796 437538 104848
rect 131114 104728 131120 104780
rect 131172 104768 131178 104780
rect 138750 104768 138756 104780
rect 131172 104740 138756 104768
rect 131172 104728 131178 104740
rect 138750 104728 138756 104740
rect 138808 104728 138814 104780
rect 411254 103504 411260 103556
rect 411312 103544 411318 103556
rect 416038 103544 416044 103556
rect 411312 103516 416044 103544
rect 411312 103504 411318 103516
rect 416038 103504 416044 103516
rect 416096 103504 416102 103556
rect 131390 103436 131396 103488
rect 131448 103476 131454 103488
rect 166258 103476 166264 103488
rect 131448 103448 166264 103476
rect 131448 103436 131454 103448
rect 166258 103436 166264 103448
rect 166316 103436 166322 103488
rect 131206 103368 131212 103420
rect 131264 103408 131270 103420
rect 145834 103408 145840 103420
rect 131264 103380 145840 103408
rect 131264 103368 131270 103380
rect 145834 103368 145840 103380
rect 145892 103368 145898 103420
rect 131114 103300 131120 103352
rect 131172 103340 131178 103352
rect 136174 103340 136180 103352
rect 131172 103312 136180 103340
rect 131172 103300 131178 103312
rect 136174 103300 136180 103312
rect 136232 103300 136238 103352
rect 435358 103028 435364 103080
rect 435416 103068 435422 103080
rect 437658 103068 437664 103080
rect 435416 103040 437664 103068
rect 435416 103028 435422 103040
rect 437658 103028 437664 103040
rect 437716 103028 437722 103080
rect 134978 102144 134984 102196
rect 135036 102184 135042 102196
rect 186314 102184 186320 102196
rect 135036 102156 186320 102184
rect 135036 102144 135042 102156
rect 186314 102144 186320 102156
rect 186372 102144 186378 102196
rect 131206 102076 131212 102128
rect 131264 102116 131270 102128
rect 138842 102116 138848 102128
rect 131264 102088 138848 102116
rect 131264 102076 131270 102088
rect 138842 102076 138848 102088
rect 138900 102076 138906 102128
rect 416130 102076 416136 102128
rect 416188 102116 416194 102128
rect 437474 102116 437480 102128
rect 416188 102088 437480 102116
rect 416188 102076 416194 102088
rect 437474 102076 437480 102088
rect 437532 102076 437538 102128
rect 134886 100716 134892 100768
rect 134944 100756 134950 100768
rect 186314 100756 186320 100768
rect 134944 100728 186320 100756
rect 134944 100716 134950 100728
rect 186314 100716 186320 100728
rect 186372 100716 186378 100768
rect 411254 100716 411260 100768
rect 411312 100756 411318 100768
rect 415118 100756 415124 100768
rect 411312 100728 415124 100756
rect 411312 100716 411318 100728
rect 415118 100716 415124 100728
rect 415176 100716 415182 100768
rect 131206 100648 131212 100700
rect 131264 100688 131270 100700
rect 164878 100688 164884 100700
rect 131264 100660 164884 100688
rect 131264 100648 131270 100660
rect 164878 100648 164884 100660
rect 164936 100648 164942 100700
rect 432598 100648 432604 100700
rect 432656 100688 432662 100700
rect 437474 100688 437480 100700
rect 432656 100660 437480 100688
rect 432656 100648 432662 100660
rect 437474 100648 437480 100660
rect 437532 100648 437538 100700
rect 540238 100648 540244 100700
rect 540296 100688 540302 100700
rect 580166 100688 580172 100700
rect 540296 100660 580172 100688
rect 540296 100648 540302 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 131114 100580 131120 100632
rect 131172 100620 131178 100632
rect 138934 100620 138940 100632
rect 131172 100592 138940 100620
rect 131172 100580 131178 100592
rect 138934 100580 138940 100592
rect 138992 100580 138998 100632
rect 140130 99424 140136 99476
rect 140188 99464 140194 99476
rect 186406 99464 186412 99476
rect 140188 99436 186412 99464
rect 140188 99424 140194 99436
rect 186406 99424 186412 99436
rect 186464 99424 186470 99476
rect 136174 99356 136180 99408
rect 136232 99396 136238 99408
rect 186314 99396 186320 99408
rect 136232 99368 186320 99396
rect 136232 99356 136238 99368
rect 186314 99356 186320 99368
rect 186372 99356 186378 99408
rect 131114 99288 131120 99340
rect 131172 99328 131178 99340
rect 162118 99328 162124 99340
rect 131172 99300 162124 99328
rect 131172 99288 131178 99300
rect 162118 99288 162124 99300
rect 162176 99288 162182 99340
rect 131206 99220 131212 99272
rect 131264 99260 131270 99272
rect 135070 99260 135076 99272
rect 131264 99232 135076 99260
rect 131264 99220 131270 99232
rect 135070 99220 135076 99232
rect 135128 99220 135134 99272
rect 133322 97996 133328 98048
rect 133380 98036 133386 98048
rect 186314 98036 186320 98048
rect 133380 98008 186320 98036
rect 133380 97996 133386 98008
rect 186314 97996 186320 98008
rect 186372 97996 186378 98048
rect 131206 97928 131212 97980
rect 131264 97968 131270 97980
rect 136266 97968 136272 97980
rect 131264 97940 136272 97968
rect 131264 97928 131270 97940
rect 136266 97928 136272 97940
rect 136324 97928 136330 97980
rect 431218 97928 431224 97980
rect 431276 97968 431282 97980
rect 437474 97968 437480 97980
rect 431276 97940 437480 97968
rect 431276 97928 431282 97940
rect 437474 97928 437480 97940
rect 437532 97928 437538 97980
rect 140222 96636 140228 96688
rect 140280 96676 140286 96688
rect 186314 96676 186320 96688
rect 140280 96648 186320 96676
rect 140280 96636 140286 96648
rect 186314 96636 186320 96648
rect 186372 96636 186378 96688
rect 131114 96568 131120 96620
rect 131172 96608 131178 96620
rect 160738 96608 160744 96620
rect 131172 96580 160744 96608
rect 131172 96568 131178 96580
rect 160738 96568 160744 96580
rect 160796 96568 160802 96620
rect 429838 96568 429844 96620
rect 429896 96608 429902 96620
rect 437474 96608 437480 96620
rect 429896 96580 437480 96608
rect 429896 96568 429902 96580
rect 437474 96568 437480 96580
rect 437532 96568 437538 96620
rect 131206 96500 131212 96552
rect 131264 96540 131270 96552
rect 139026 96540 139032 96552
rect 131264 96512 139032 96540
rect 131264 96500 131270 96512
rect 139026 96500 139032 96512
rect 139084 96500 139090 96552
rect 131390 95888 131396 95940
rect 131448 95928 131454 95940
rect 133782 95928 133788 95940
rect 131448 95900 133788 95928
rect 131448 95888 131454 95900
rect 133782 95888 133788 95900
rect 133840 95888 133846 95940
rect 411254 95820 411260 95872
rect 411312 95860 411318 95872
rect 415210 95860 415216 95872
rect 411312 95832 415216 95860
rect 411312 95820 411318 95832
rect 415210 95820 415216 95832
rect 415268 95820 415274 95872
rect 144730 95208 144736 95260
rect 144788 95248 144794 95260
rect 186314 95248 186320 95260
rect 144788 95220 186320 95248
rect 144788 95208 144794 95220
rect 186314 95208 186320 95220
rect 186372 95208 186378 95260
rect 131114 95140 131120 95192
rect 131172 95180 131178 95192
rect 145926 95180 145932 95192
rect 131172 95152 145932 95180
rect 131172 95140 131178 95152
rect 145926 95140 145932 95152
rect 145984 95140 145990 95192
rect 428458 95140 428464 95192
rect 428516 95180 428522 95192
rect 437474 95180 437480 95192
rect 428516 95152 437480 95180
rect 428516 95140 428522 95152
rect 437474 95140 437480 95152
rect 437532 95140 437538 95192
rect 131206 95072 131212 95124
rect 131264 95112 131270 95124
rect 137462 95112 137468 95124
rect 131264 95084 137468 95112
rect 131264 95072 131270 95084
rect 137462 95072 137468 95084
rect 137520 95072 137526 95124
rect 411254 93916 411260 93968
rect 411312 93956 411318 93968
rect 413370 93956 413376 93968
rect 411312 93928 413376 93956
rect 411312 93916 411318 93928
rect 413370 93916 413376 93928
rect 413428 93916 413434 93968
rect 133506 93848 133512 93900
rect 133564 93888 133570 93900
rect 186314 93888 186320 93900
rect 133564 93860 186320 93888
rect 133564 93848 133570 93860
rect 186314 93848 186320 93860
rect 186372 93848 186378 93900
rect 131206 93780 131212 93832
rect 131264 93820 131270 93832
rect 147122 93820 147128 93832
rect 131264 93792 147128 93820
rect 131264 93780 131270 93792
rect 147122 93780 147128 93792
rect 147180 93780 147186 93832
rect 425698 93780 425704 93832
rect 425756 93820 425762 93832
rect 437474 93820 437480 93832
rect 425756 93792 437480 93820
rect 425756 93780 425762 93792
rect 437474 93780 437480 93792
rect 437532 93780 437538 93832
rect 131114 93712 131120 93764
rect 131172 93752 131178 93764
rect 146018 93752 146024 93764
rect 131172 93724 146024 93752
rect 131172 93712 131178 93724
rect 146018 93712 146024 93724
rect 146076 93712 146082 93764
rect 138658 92556 138664 92608
rect 138716 92596 138722 92608
rect 186406 92596 186412 92608
rect 138716 92568 186412 92596
rect 138716 92556 138722 92568
rect 186406 92556 186412 92568
rect 186464 92556 186470 92608
rect 131942 92488 131948 92540
rect 132000 92528 132006 92540
rect 186314 92528 186320 92540
rect 132000 92500 186320 92528
rect 132000 92488 132006 92500
rect 186314 92488 186320 92500
rect 186372 92488 186378 92540
rect 131114 92420 131120 92472
rect 131172 92460 131178 92472
rect 144178 92460 144184 92472
rect 131172 92432 144184 92460
rect 131172 92420 131178 92432
rect 144178 92420 144184 92432
rect 144236 92420 144242 92472
rect 411254 92420 411260 92472
rect 411312 92460 411318 92472
rect 419350 92460 419356 92472
rect 411312 92432 419356 92460
rect 411312 92420 411318 92432
rect 419350 92420 419356 92432
rect 419408 92420 419414 92472
rect 424318 92420 424324 92472
rect 424376 92460 424382 92472
rect 437474 92460 437480 92472
rect 424376 92432 437480 92460
rect 424376 92420 424382 92432
rect 437474 92420 437480 92432
rect 437532 92420 437538 92472
rect 131206 92352 131212 92404
rect 131264 92392 131270 92404
rect 137554 92392 137560 92404
rect 131264 92364 137560 92392
rect 131264 92352 131270 92364
rect 137554 92352 137560 92364
rect 137612 92352 137618 92404
rect 133414 91060 133420 91112
rect 133472 91100 133478 91112
rect 186314 91100 186320 91112
rect 133472 91072 186320 91100
rect 133472 91060 133478 91072
rect 186314 91060 186320 91072
rect 186372 91060 186378 91112
rect 132218 90992 132224 91044
rect 132276 91032 132282 91044
rect 144270 91032 144276 91044
rect 132276 91004 144276 91032
rect 132276 90992 132282 91004
rect 144270 90992 144276 91004
rect 144328 90992 144334 91044
rect 421742 90992 421748 91044
rect 421800 91032 421806 91044
rect 437474 91032 437480 91044
rect 421800 91004 437480 91032
rect 421800 90992 421806 91004
rect 437474 90992 437480 91004
rect 437532 90992 437538 91044
rect 131206 90924 131212 90976
rect 131264 90964 131270 90976
rect 143074 90964 143080 90976
rect 131264 90936 143080 90964
rect 131264 90924 131270 90936
rect 143074 90924 143080 90936
rect 143132 90924 143138 90976
rect 411254 89768 411260 89820
rect 411312 89808 411318 89820
rect 413370 89808 413376 89820
rect 411312 89780 413376 89808
rect 411312 89768 411318 89780
rect 413370 89768 413376 89780
rect 413428 89768 413434 89820
rect 138750 89700 138756 89752
rect 138808 89740 138814 89752
rect 186314 89740 186320 89752
rect 138808 89712 186320 89740
rect 138808 89700 138814 89712
rect 186314 89700 186320 89712
rect 186372 89700 186378 89752
rect 131114 89632 131120 89684
rect 131172 89672 131178 89684
rect 144362 89672 144368 89684
rect 131172 89644 144368 89672
rect 131172 89632 131178 89644
rect 144362 89632 144368 89644
rect 144420 89632 144426 89684
rect 418982 89632 418988 89684
rect 419040 89672 419046 89684
rect 437474 89672 437480 89684
rect 419040 89644 437480 89672
rect 419040 89632 419046 89644
rect 437474 89632 437480 89644
rect 437532 89632 437538 89684
rect 131206 89564 131212 89616
rect 131264 89604 131270 89616
rect 141602 89604 141608 89616
rect 131264 89576 141608 89604
rect 131264 89564 131270 89576
rect 141602 89564 141608 89576
rect 141660 89564 141666 89616
rect 132126 88340 132132 88392
rect 132184 88380 132190 88392
rect 186314 88380 186320 88392
rect 132184 88352 186320 88380
rect 132184 88340 132190 88352
rect 186314 88340 186320 88352
rect 186372 88340 186378 88392
rect 131114 88272 131120 88324
rect 131172 88312 131178 88324
rect 187326 88312 187332 88324
rect 131172 88284 187332 88312
rect 131172 88272 131178 88284
rect 187326 88272 187332 88284
rect 187384 88272 187390 88324
rect 411254 88272 411260 88324
rect 411312 88312 411318 88324
rect 419258 88312 419264 88324
rect 411312 88284 419264 88312
rect 411312 88272 411318 88284
rect 419258 88272 419264 88284
rect 419316 88272 419322 88324
rect 420270 88272 420276 88324
rect 420328 88312 420334 88324
rect 437474 88312 437480 88324
rect 420328 88284 437480 88312
rect 420328 88272 420334 88284
rect 437474 88272 437480 88284
rect 437532 88272 437538 88324
rect 131206 88204 131212 88256
rect 131264 88244 131270 88256
rect 142982 88244 142988 88256
rect 131264 88216 142988 88244
rect 131264 88204 131270 88216
rect 142982 88204 142988 88216
rect 143040 88204 143046 88256
rect 131298 88136 131304 88188
rect 131356 88176 131362 88188
rect 137646 88176 137652 88188
rect 131356 88148 137652 88176
rect 131356 88136 131362 88148
rect 137646 88136 137652 88148
rect 137704 88136 137710 88188
rect 133598 86980 133604 87032
rect 133656 87020 133662 87032
rect 186314 87020 186320 87032
rect 133656 86992 186320 87020
rect 133656 86980 133662 86992
rect 186314 86980 186320 86992
rect 186372 86980 186378 87032
rect 131114 86912 131120 86964
rect 131172 86952 131178 86964
rect 143166 86952 143172 86964
rect 131172 86924 143172 86952
rect 131172 86912 131178 86924
rect 143166 86912 143172 86924
rect 143224 86912 143230 86964
rect 131206 86844 131212 86896
rect 131264 86884 131270 86896
rect 141694 86884 141700 86896
rect 131264 86856 141700 86884
rect 131264 86844 131270 86856
rect 141694 86844 141700 86856
rect 141752 86844 141758 86896
rect 411254 86436 411260 86488
rect 411312 86476 411318 86488
rect 413830 86476 413836 86488
rect 411312 86448 413836 86476
rect 411312 86436 411318 86448
rect 413830 86436 413836 86448
rect 413888 86436 413894 86488
rect 131666 85552 131672 85604
rect 131724 85592 131730 85604
rect 186314 85592 186320 85604
rect 131724 85564 186320 85592
rect 131724 85552 131730 85564
rect 186314 85552 186320 85564
rect 186372 85552 186378 85604
rect 131114 85484 131120 85536
rect 131172 85524 131178 85536
rect 143258 85524 143264 85536
rect 131172 85496 143264 85524
rect 131172 85484 131178 85496
rect 143258 85484 143264 85496
rect 143316 85484 143322 85536
rect 417418 85484 417424 85536
rect 417476 85524 417482 85536
rect 437474 85524 437480 85536
rect 417476 85496 437480 85524
rect 417476 85484 417482 85496
rect 437474 85484 437480 85496
rect 437532 85484 437538 85536
rect 131206 85416 131212 85468
rect 131264 85456 131270 85468
rect 137738 85456 137744 85468
rect 131264 85428 137744 85456
rect 131264 85416 131270 85428
rect 137738 85416 137744 85428
rect 137796 85416 137802 85468
rect 142982 84192 142988 84244
rect 143040 84232 143046 84244
rect 186314 84232 186320 84244
rect 143040 84204 186320 84232
rect 143040 84192 143046 84204
rect 186314 84192 186320 84204
rect 186372 84192 186378 84244
rect 131114 84124 131120 84176
rect 131172 84164 131178 84176
rect 141878 84164 141884 84176
rect 131172 84136 141884 84164
rect 131172 84124 131178 84136
rect 141878 84124 141884 84136
rect 141936 84124 141942 84176
rect 411254 84124 411260 84176
rect 411312 84164 411318 84176
rect 413738 84164 413744 84176
rect 411312 84136 413744 84164
rect 411312 84124 411318 84136
rect 413738 84124 413744 84136
rect 413796 84124 413802 84176
rect 420178 84124 420184 84176
rect 420236 84164 420242 84176
rect 437474 84164 437480 84176
rect 420236 84136 437480 84164
rect 420236 84124 420242 84136
rect 437474 84124 437480 84136
rect 437532 84124 437538 84176
rect 131206 84056 131212 84108
rect 131264 84096 131270 84108
rect 140406 84096 140412 84108
rect 131264 84068 140412 84096
rect 131264 84056 131270 84068
rect 140406 84056 140412 84068
rect 140464 84056 140470 84108
rect 131574 83988 131580 84040
rect 131632 84028 131638 84040
rect 137830 84028 137836 84040
rect 131632 84000 137836 84028
rect 131632 83988 131638 84000
rect 137830 83988 137836 84000
rect 137888 83988 137894 84040
rect 131206 82764 131212 82816
rect 131264 82804 131270 82816
rect 187418 82804 187424 82816
rect 131264 82776 187424 82804
rect 131264 82764 131270 82776
rect 187418 82764 187424 82776
rect 187476 82764 187482 82816
rect 417602 82764 417608 82816
rect 417660 82804 417666 82816
rect 437474 82804 437480 82816
rect 417660 82776 437480 82804
rect 417660 82764 417666 82776
rect 437474 82764 437480 82776
rect 437532 82764 437538 82816
rect 131114 82696 131120 82748
rect 131172 82736 131178 82748
rect 144454 82736 144460 82748
rect 131172 82708 144460 82736
rect 131172 82696 131178 82708
rect 144454 82696 144460 82708
rect 144512 82696 144518 82748
rect 132218 81404 132224 81456
rect 132276 81444 132282 81456
rect 186314 81444 186320 81456
rect 132276 81416 186320 81444
rect 132276 81404 132282 81416
rect 186314 81404 186320 81416
rect 186372 81404 186378 81456
rect 411254 81404 411260 81456
rect 411312 81444 411318 81456
rect 439498 81444 439504 81456
rect 411312 81416 439504 81444
rect 411312 81404 411318 81416
rect 439498 81404 439504 81416
rect 439556 81404 439562 81456
rect 131206 81336 131212 81388
rect 131264 81376 131270 81388
rect 141786 81376 141792 81388
rect 131264 81348 141792 81376
rect 131264 81336 131270 81348
rect 141786 81336 141792 81348
rect 141844 81336 141850 81388
rect 420362 81336 420368 81388
rect 420420 81376 420426 81388
rect 437474 81376 437480 81388
rect 420420 81348 437480 81376
rect 420420 81336 420426 81348
rect 437474 81336 437480 81348
rect 437532 81336 437538 81388
rect 131114 81268 131120 81320
rect 131172 81308 131178 81320
rect 140498 81308 140504 81320
rect 131172 81280 140504 81308
rect 131172 81268 131178 81280
rect 140498 81268 140504 81280
rect 140556 81268 140562 81320
rect 133690 80044 133696 80096
rect 133748 80084 133754 80096
rect 186314 80084 186320 80096
rect 133748 80056 186320 80084
rect 133748 80044 133754 80056
rect 186314 80044 186320 80056
rect 186372 80044 186378 80096
rect 131298 79976 131304 80028
rect 131356 80016 131362 80028
rect 187510 80016 187516 80028
rect 131356 79988 187516 80016
rect 131356 79976 131362 79988
rect 187510 79976 187516 79988
rect 187568 79976 187574 80028
rect 417510 79976 417516 80028
rect 417568 80016 417574 80028
rect 437474 80016 437480 80028
rect 417568 79988 437480 80016
rect 417568 79976 417574 79988
rect 437474 79976 437480 79988
rect 437532 79976 437538 80028
rect 131206 79908 131212 79960
rect 131264 79948 131270 79960
rect 144546 79948 144552 79960
rect 131264 79920 144552 79948
rect 131264 79908 131270 79920
rect 144546 79908 144552 79920
rect 144604 79908 144610 79960
rect 131114 79840 131120 79892
rect 131172 79880 131178 79892
rect 141970 79880 141976 79892
rect 131172 79852 141976 79880
rect 131172 79840 131178 79852
rect 141970 79840 141976 79852
rect 142028 79840 142034 79892
rect 131666 79296 131672 79348
rect 131724 79336 131730 79348
rect 132034 79336 132040 79348
rect 131724 79308 132040 79336
rect 131724 79296 131730 79308
rect 132034 79296 132040 79308
rect 132092 79296 132098 79348
rect 135070 78684 135076 78736
rect 135128 78724 135134 78736
rect 186314 78724 186320 78736
rect 135128 78696 186320 78724
rect 135128 78684 135134 78696
rect 186314 78684 186320 78696
rect 186372 78684 186378 78736
rect 131206 78616 131212 78668
rect 131264 78656 131270 78668
rect 144638 78656 144644 78668
rect 131264 78628 144644 78656
rect 131264 78616 131270 78628
rect 144638 78616 144644 78628
rect 144696 78616 144702 78668
rect 419074 78616 419080 78668
rect 419132 78656 419138 78668
rect 437474 78656 437480 78668
rect 419132 78628 437480 78656
rect 419132 78616 419138 78628
rect 437474 78616 437480 78628
rect 437532 78616 437538 78668
rect 131114 78548 131120 78600
rect 131172 78588 131178 78600
rect 141418 78588 141424 78600
rect 131172 78560 141424 78588
rect 131172 78548 131178 78560
rect 141418 78548 141424 78560
rect 141476 78548 141482 78600
rect 411254 78208 411260 78260
rect 411312 78248 411318 78260
rect 413646 78248 413652 78260
rect 411312 78220 413652 78248
rect 411312 78208 411318 78220
rect 413646 78208 413652 78220
rect 413704 78208 413710 78260
rect 141510 77256 141516 77308
rect 141568 77296 141574 77308
rect 186314 77296 186320 77308
rect 141568 77268 186320 77296
rect 141568 77256 141574 77268
rect 186314 77256 186320 77268
rect 186372 77256 186378 77308
rect 417694 77188 417700 77240
rect 417752 77228 417758 77240
rect 437474 77228 437480 77240
rect 417752 77200 437480 77228
rect 417752 77188 417758 77200
rect 437474 77188 437480 77200
rect 437532 77188 437538 77240
rect 131298 77120 131304 77172
rect 131356 77160 131362 77172
rect 142798 77160 142804 77172
rect 131356 77132 142804 77160
rect 131356 77120 131362 77132
rect 142798 77120 142804 77132
rect 142856 77120 142862 77172
rect 131206 77052 131212 77104
rect 131264 77092 131270 77104
rect 186958 77092 186964 77104
rect 131264 77064 186964 77092
rect 131264 77052 131270 77064
rect 186958 77052 186964 77064
rect 187016 77052 187022 77104
rect 411254 76712 411260 76764
rect 411312 76752 411318 76764
rect 413462 76752 413468 76764
rect 411312 76724 413468 76752
rect 411312 76712 411318 76724
rect 413462 76712 413468 76724
rect 413520 76712 413526 76764
rect 131666 76576 131672 76628
rect 131724 76616 131730 76628
rect 134610 76616 134616 76628
rect 131724 76588 134616 76616
rect 131724 76576 131730 76588
rect 134610 76576 134616 76588
rect 134668 76576 134674 76628
rect 131206 75828 131212 75880
rect 131264 75868 131270 75880
rect 142890 75868 142896 75880
rect 131264 75840 142896 75868
rect 131264 75828 131270 75840
rect 142890 75828 142896 75840
rect 142948 75828 142954 75880
rect 134610 74604 134616 74656
rect 134668 74644 134674 74656
rect 186406 74644 186412 74656
rect 134668 74616 186412 74644
rect 134668 74604 134674 74616
rect 186406 74604 186412 74616
rect 186464 74604 186470 74656
rect 133782 74536 133788 74588
rect 133840 74576 133846 74588
rect 186314 74576 186320 74588
rect 133840 74548 186320 74576
rect 133840 74536 133846 74548
rect 186314 74536 186320 74548
rect 186372 74536 186378 74588
rect 131850 74468 131856 74520
rect 131908 74508 131914 74520
rect 134518 74508 134524 74520
rect 131908 74480 134524 74508
rect 131908 74468 131914 74480
rect 134518 74468 134524 74480
rect 134576 74468 134582 74520
rect 414934 74468 414940 74520
rect 414992 74508 414998 74520
rect 437474 74508 437480 74520
rect 414992 74480 437480 74508
rect 414992 74468 414998 74480
rect 437474 74468 437480 74480
rect 437532 74468 437538 74520
rect 411254 74196 411260 74248
rect 411312 74236 411318 74248
rect 413554 74236 413560 74248
rect 411312 74208 413560 74236
rect 411312 74196 411318 74208
rect 413554 74196 413560 74208
rect 413612 74196 413618 74248
rect 131298 73108 131304 73160
rect 131356 73148 131362 73160
rect 187050 73148 187056 73160
rect 131356 73120 187056 73148
rect 131356 73108 131362 73120
rect 187050 73108 187056 73120
rect 187108 73108 187114 73160
rect 411254 73108 411260 73160
rect 411312 73148 411318 73160
rect 438486 73148 438492 73160
rect 411312 73120 438492 73148
rect 411312 73108 411318 73120
rect 438486 73108 438492 73120
rect 438544 73108 438550 73160
rect 131206 73040 131212 73092
rect 131264 73080 131270 73092
rect 135898 73080 135904 73092
rect 131264 73052 135904 73080
rect 131264 73040 131270 73052
rect 135898 73040 135904 73052
rect 135956 73040 135962 73092
rect 417786 73040 417792 73092
rect 417844 73080 417850 73092
rect 437474 73080 437480 73092
rect 417844 73052 437480 73080
rect 417844 73040 417850 73052
rect 437474 73040 437480 73052
rect 437532 73040 437538 73092
rect 131114 72972 131120 73024
rect 131172 73012 131178 73024
rect 134702 73012 134708 73024
rect 131172 72984 134708 73012
rect 131172 72972 131178 72984
rect 134702 72972 134708 72984
rect 134760 72972 134766 73024
rect 151078 71748 151084 71800
rect 151136 71788 151142 71800
rect 186314 71788 186320 71800
rect 151136 71760 186320 71788
rect 151136 71748 151142 71760
rect 186314 71748 186320 71760
rect 186372 71748 186378 71800
rect 131114 71680 131120 71732
rect 131172 71720 131178 71732
rect 133230 71720 133236 71732
rect 131172 71692 133236 71720
rect 131172 71680 131178 71692
rect 133230 71680 133236 71692
rect 133288 71680 133294 71732
rect 415026 71680 415032 71732
rect 415084 71720 415090 71732
rect 437474 71720 437480 71732
rect 415084 71692 437480 71720
rect 415084 71680 415090 71692
rect 437474 71680 437480 71692
rect 437532 71680 437538 71732
rect 131206 71612 131212 71664
rect 131264 71652 131270 71664
rect 135990 71652 135996 71664
rect 131264 71624 135996 71652
rect 131264 71612 131270 71624
rect 135990 71612 135996 71624
rect 136048 71612 136054 71664
rect 134518 70388 134524 70440
rect 134576 70428 134582 70440
rect 186314 70428 186320 70440
rect 134576 70400 186320 70428
rect 134576 70388 134582 70400
rect 186314 70388 186320 70400
rect 186372 70388 186378 70440
rect 131206 70320 131212 70372
rect 131264 70360 131270 70372
rect 140038 70360 140044 70372
rect 131264 70332 140044 70360
rect 131264 70320 131270 70332
rect 140038 70320 140044 70332
rect 140096 70320 140102 70372
rect 421834 70320 421840 70372
rect 421892 70360 421898 70372
rect 437474 70360 437480 70372
rect 421892 70332 437480 70360
rect 421892 70320 421898 70332
rect 437474 70320 437480 70332
rect 437532 70320 437538 70372
rect 131114 70252 131120 70304
rect 131172 70292 131178 70304
rect 136082 70292 136088 70304
rect 131172 70264 136088 70292
rect 131172 70252 131178 70264
rect 136082 70252 136088 70264
rect 136140 70252 136146 70304
rect 131574 69640 131580 69692
rect 131632 69680 131638 69692
rect 132034 69680 132040 69692
rect 131632 69652 132040 69680
rect 131632 69640 131638 69652
rect 132034 69640 132040 69652
rect 132092 69640 132098 69692
rect 137278 69096 137284 69148
rect 137336 69136 137342 69148
rect 186314 69136 186320 69148
rect 137336 69108 186320 69136
rect 137336 69096 137342 69108
rect 186314 69096 186320 69108
rect 186372 69096 186378 69148
rect 131850 69028 131856 69080
rect 131908 69068 131914 69080
rect 186406 69068 186412 69080
rect 131908 69040 186412 69068
rect 131908 69028 131914 69040
rect 186406 69028 186412 69040
rect 186464 69028 186470 69080
rect 411346 69028 411352 69080
rect 411404 69068 411410 69080
rect 418982 69068 418988 69080
rect 411404 69040 418988 69068
rect 411404 69028 411410 69040
rect 418982 69028 418988 69040
rect 419040 69028 419046 69080
rect 131390 68960 131396 69012
rect 131448 69000 131454 69012
rect 187142 69000 187148 69012
rect 131448 68972 187148 69000
rect 131448 68960 131454 68972
rect 187142 68960 187148 68972
rect 187200 68960 187206 69012
rect 411254 68960 411260 69012
rect 411312 69000 411318 69012
rect 438394 69000 438400 69012
rect 411312 68972 438400 69000
rect 411312 68960 411318 68972
rect 438394 68960 438400 68972
rect 438452 68960 438458 69012
rect 131206 68892 131212 68944
rect 131264 68932 131270 68944
rect 134794 68932 134800 68944
rect 131264 68904 134800 68932
rect 131264 68892 131270 68904
rect 134794 68892 134800 68904
rect 134852 68892 134858 68944
rect 417878 68892 417884 68944
rect 417936 68932 417942 68944
rect 437474 68932 437480 68944
rect 417936 68904 437480 68932
rect 417936 68892 417942 68904
rect 437474 68892 437480 68904
rect 437532 68892 437538 68944
rect 131114 68824 131120 68876
rect 131172 68864 131178 68876
rect 134978 68864 134984 68876
rect 131172 68836 134984 68864
rect 131172 68824 131178 68836
rect 134978 68824 134984 68836
rect 135036 68824 135042 68876
rect 148318 67600 148324 67652
rect 148376 67640 148382 67652
rect 186314 67640 186320 67652
rect 148376 67612 186320 67640
rect 148376 67600 148382 67612
rect 186314 67600 186320 67612
rect 186372 67600 186378 67652
rect 131114 67532 131120 67584
rect 131172 67572 131178 67584
rect 140130 67572 140136 67584
rect 131172 67544 140136 67572
rect 131172 67532 131178 67544
rect 140130 67532 140136 67544
rect 140188 67532 140194 67584
rect 429930 67532 429936 67584
rect 429988 67572 429994 67584
rect 437474 67572 437480 67584
rect 429988 67544 437480 67572
rect 429988 67532 429994 67544
rect 437474 67532 437480 67544
rect 437532 67532 437538 67584
rect 131206 67328 131212 67380
rect 131264 67368 131270 67380
rect 134886 67368 134892 67380
rect 131264 67340 134892 67368
rect 131264 67328 131270 67340
rect 134886 67328 134892 67340
rect 134944 67328 134950 67380
rect 133230 66240 133236 66292
rect 133288 66280 133294 66292
rect 186314 66280 186320 66292
rect 133288 66252 186320 66280
rect 133288 66240 133294 66252
rect 186314 66240 186320 66252
rect 186372 66240 186378 66292
rect 411254 66240 411260 66292
rect 411312 66280 411318 66292
rect 436738 66280 436744 66292
rect 411312 66252 436744 66280
rect 411312 66240 411318 66252
rect 436738 66240 436744 66252
rect 436796 66240 436802 66292
rect 131206 66172 131212 66224
rect 131264 66212 131270 66224
rect 136174 66212 136180 66224
rect 131264 66184 136180 66212
rect 131264 66172 131270 66184
rect 136174 66172 136180 66184
rect 136232 66172 136238 66224
rect 421926 66172 421932 66224
rect 421984 66212 421990 66224
rect 437474 66212 437480 66224
rect 421984 66184 437480 66212
rect 421984 66172 421990 66184
rect 437474 66172 437480 66184
rect 437532 66172 437538 66224
rect 131114 66104 131120 66156
rect 131172 66144 131178 66156
rect 133322 66144 133328 66156
rect 131172 66116 133328 66144
rect 131172 66104 131178 66116
rect 133322 66104 133328 66116
rect 133380 66104 133386 66156
rect 132126 64880 132132 64932
rect 132184 64920 132190 64932
rect 186314 64920 186320 64932
rect 132184 64892 186320 64920
rect 132184 64880 132190 64892
rect 186314 64880 186320 64892
rect 186372 64880 186378 64932
rect 131298 64812 131304 64864
rect 131356 64852 131362 64864
rect 144730 64852 144736 64864
rect 131356 64824 144736 64852
rect 131356 64812 131362 64824
rect 144730 64812 144736 64824
rect 144788 64812 144794 64864
rect 431310 64812 431316 64864
rect 431368 64852 431374 64864
rect 437474 64852 437480 64864
rect 431368 64824 437480 64852
rect 431368 64812 431374 64824
rect 437474 64812 437480 64824
rect 437532 64812 437538 64864
rect 131206 64744 131212 64796
rect 131264 64784 131270 64796
rect 140222 64784 140228 64796
rect 131264 64756 140228 64784
rect 131264 64744 131270 64756
rect 140222 64744 140228 64756
rect 140280 64744 140286 64796
rect 131114 64676 131120 64728
rect 131172 64716 131178 64728
rect 133506 64716 133512 64728
rect 131172 64688 133512 64716
rect 131172 64676 131178 64688
rect 133506 64676 133512 64688
rect 133564 64676 133570 64728
rect 411254 64472 411260 64524
rect 411312 64512 411318 64524
rect 413278 64512 413284 64524
rect 411312 64484 413284 64512
rect 411312 64472 411318 64484
rect 413278 64472 413284 64484
rect 413336 64472 413342 64524
rect 146938 63520 146944 63572
rect 146996 63560 147002 63572
rect 186314 63560 186320 63572
rect 146996 63532 186320 63560
rect 146996 63520 147002 63532
rect 186314 63520 186320 63532
rect 186372 63520 186378 63572
rect 131206 63452 131212 63504
rect 131264 63492 131270 63504
rect 138658 63492 138664 63504
rect 131264 63464 138664 63492
rect 131264 63452 131270 63464
rect 138658 63452 138664 63464
rect 138716 63452 138722 63504
rect 411254 63452 411260 63504
rect 411312 63492 411318 63504
rect 438302 63492 438308 63504
rect 411312 63464 438308 63492
rect 411312 63452 411318 63464
rect 438302 63452 438308 63464
rect 438360 63452 438366 63504
rect 132402 62092 132408 62144
rect 132460 62132 132466 62144
rect 186314 62132 186320 62144
rect 132460 62104 186320 62132
rect 132460 62092 132466 62104
rect 186314 62092 186320 62104
rect 186372 62092 186378 62144
rect 131114 62024 131120 62076
rect 131172 62064 131178 62076
rect 138750 62064 138756 62076
rect 131172 62036 138756 62064
rect 131172 62024 131178 62036
rect 138750 62024 138756 62036
rect 138808 62024 138814 62076
rect 422018 62024 422024 62076
rect 422076 62064 422082 62076
rect 437474 62064 437480 62076
rect 422076 62036 437480 62064
rect 422076 62024 422082 62036
rect 437474 62024 437480 62036
rect 437532 62024 437538 62076
rect 131206 61956 131212 62008
rect 131264 61996 131270 62008
rect 133414 61996 133420 62008
rect 131264 61968 133420 61996
rect 131264 61956 131270 61968
rect 133414 61956 133420 61968
rect 133472 61956 133478 62008
rect 144178 60732 144184 60784
rect 144236 60772 144242 60784
rect 186314 60772 186320 60784
rect 144236 60744 186320 60772
rect 144236 60732 144242 60744
rect 186314 60732 186320 60744
rect 186372 60732 186378 60784
rect 131114 60664 131120 60716
rect 131172 60704 131178 60716
rect 187234 60704 187240 60716
rect 131172 60676 187240 60704
rect 131172 60664 131178 60676
rect 187234 60664 187240 60676
rect 187292 60664 187298 60716
rect 432690 60664 432696 60716
rect 432748 60704 432754 60716
rect 437474 60704 437480 60716
rect 432748 60676 437480 60704
rect 432748 60664 432754 60676
rect 437474 60664 437480 60676
rect 437532 60664 437538 60716
rect 544378 60664 544384 60716
rect 544436 60704 544442 60716
rect 579798 60704 579804 60716
rect 544436 60676 579804 60704
rect 544436 60664 544442 60676
rect 579798 60664 579804 60676
rect 579856 60664 579862 60716
rect 131206 60596 131212 60648
rect 131264 60636 131270 60648
rect 133598 60636 133604 60648
rect 131264 60608 133604 60636
rect 131264 60596 131270 60608
rect 133598 60596 133604 60608
rect 133656 60596 133662 60648
rect 411254 59372 411260 59424
rect 411312 59412 411318 59424
rect 417418 59412 417424 59424
rect 411312 59384 417424 59412
rect 411312 59372 411318 59384
rect 417418 59372 417424 59384
rect 417476 59372 417482 59424
rect 131206 59304 131212 59356
rect 131264 59344 131270 59356
rect 142982 59344 142988 59356
rect 131264 59316 142988 59344
rect 131264 59304 131270 59316
rect 142982 59304 142988 59316
rect 143040 59304 143046 59356
rect 420454 59304 420460 59356
rect 420512 59344 420518 59356
rect 437474 59344 437480 59356
rect 420512 59316 437480 59344
rect 420512 59304 420518 59316
rect 437474 59304 437480 59316
rect 437532 59304 437538 59356
rect 131942 57944 131948 57996
rect 132000 57984 132006 57996
rect 186314 57984 186320 57996
rect 132000 57956 186320 57984
rect 132000 57944 132006 57956
rect 186314 57944 186320 57956
rect 186372 57944 186378 57996
rect 411254 57944 411260 57996
rect 411312 57984 411318 57996
rect 439590 57984 439596 57996
rect 411312 57956 439596 57984
rect 411312 57944 411318 57956
rect 439590 57944 439596 57956
rect 439648 57944 439654 57996
rect 131206 57876 131212 57928
rect 131264 57916 131270 57928
rect 187326 57916 187332 57928
rect 131264 57888 187332 57916
rect 131264 57876 131270 57888
rect 187326 57876 187332 57888
rect 187384 57876 187390 57928
rect 412174 57876 412180 57928
rect 412232 57916 412238 57928
rect 437474 57916 437480 57928
rect 412232 57888 437480 57916
rect 412232 57876 412238 57888
rect 437474 57876 437480 57888
rect 437532 57876 437538 57928
rect 131206 57332 131212 57384
rect 131264 57372 131270 57384
rect 133690 57372 133696 57384
rect 131264 57344 133696 57372
rect 131264 57332 131270 57344
rect 133690 57332 133696 57344
rect 133748 57332 133754 57384
rect 133322 56584 133328 56636
rect 133380 56624 133386 56636
rect 186314 56624 186320 56636
rect 133380 56596 186320 56624
rect 133380 56584 133386 56596
rect 186314 56584 186320 56596
rect 186372 56584 186378 56636
rect 131206 56516 131212 56568
rect 131264 56556 131270 56568
rect 187418 56556 187424 56568
rect 131264 56528 187424 56556
rect 131264 56516 131270 56528
rect 187418 56516 187424 56528
rect 187476 56516 187482 56568
rect 420546 56516 420552 56568
rect 420604 56556 420610 56568
rect 437474 56556 437480 56568
rect 420604 56528 437480 56556
rect 420604 56516 420610 56528
rect 437474 56516 437480 56528
rect 437532 56516 437538 56568
rect 131114 56448 131120 56500
rect 131172 56488 131178 56500
rect 135070 56488 135076 56500
rect 131172 56460 135076 56488
rect 131172 56448 131178 56460
rect 135070 56448 135076 56460
rect 135128 56448 135134 56500
rect 132034 55224 132040 55276
rect 132092 55264 132098 55276
rect 186314 55264 186320 55276
rect 132092 55236 186320 55264
rect 132092 55224 132098 55236
rect 186314 55224 186320 55236
rect 186372 55224 186378 55276
rect 131206 55156 131212 55208
rect 131264 55196 131270 55208
rect 187510 55196 187516 55208
rect 131264 55168 187516 55196
rect 131264 55156 131270 55168
rect 187510 55156 187516 55168
rect 187568 55156 187574 55208
rect 132126 55088 132132 55140
rect 132184 55128 132190 55140
rect 141510 55128 141516 55140
rect 132184 55100 141516 55128
rect 132184 55088 132190 55100
rect 141510 55088 141516 55100
rect 141568 55088 141574 55140
rect 435450 54680 435456 54732
rect 435508 54720 435514 54732
rect 437750 54720 437756 54732
rect 435508 54692 437756 54720
rect 435508 54680 435514 54692
rect 437750 54680 437756 54692
rect 437808 54680 437814 54732
rect 411254 54000 411260 54052
rect 411312 54040 411318 54052
rect 413462 54040 413468 54052
rect 411312 54012 413468 54040
rect 411312 54000 411318 54012
rect 413462 54000 413468 54012
rect 413520 54000 413526 54052
rect 133414 53796 133420 53848
rect 133472 53836 133478 53848
rect 186314 53836 186320 53848
rect 133472 53808 186320 53836
rect 133472 53796 133478 53808
rect 186314 53796 186320 53808
rect 186372 53796 186378 53848
rect 131666 53728 131672 53780
rect 131724 53768 131730 53780
rect 133782 53768 133788 53780
rect 131724 53740 133788 53768
rect 131724 53728 131730 53740
rect 133782 53728 133788 53740
rect 133840 53728 133846 53780
rect 416222 53728 416228 53780
rect 416280 53768 416286 53780
rect 437474 53768 437480 53780
rect 416280 53740 437480 53768
rect 416280 53728 416286 53740
rect 437474 53728 437480 53740
rect 437532 53728 437538 53780
rect 131206 53660 131212 53712
rect 131264 53700 131270 53712
rect 134610 53700 134616 53712
rect 131264 53672 134616 53700
rect 131264 53660 131270 53672
rect 134610 53660 134616 53672
rect 134668 53660 134674 53712
rect 131114 53592 131120 53644
rect 131172 53632 131178 53644
rect 186958 53632 186964 53644
rect 131172 53604 186964 53632
rect 131172 53592 131178 53604
rect 186958 53592 186964 53604
rect 187016 53592 187022 53644
rect 411254 52504 411260 52556
rect 411312 52544 411318 52556
rect 413278 52544 413284 52556
rect 411312 52516 413284 52544
rect 411312 52504 411318 52516
rect 413278 52504 413284 52516
rect 413336 52504 413342 52556
rect 132218 52368 132224 52420
rect 132276 52408 132282 52420
rect 151078 52408 151084 52420
rect 132276 52380 151084 52408
rect 132276 52368 132282 52380
rect 151078 52368 151084 52380
rect 151136 52368 151142 52420
rect 428550 52368 428556 52420
rect 428608 52408 428614 52420
rect 437474 52408 437480 52420
rect 428608 52380 437480 52408
rect 428608 52368 428614 52380
rect 437474 52368 437480 52380
rect 437532 52368 437538 52420
rect 131206 52300 131212 52352
rect 131264 52340 131270 52352
rect 134518 52340 134524 52352
rect 131264 52312 134524 52340
rect 131264 52300 131270 52312
rect 134518 52300 134524 52312
rect 134576 52300 134582 52352
rect 132218 51076 132224 51128
rect 132276 51116 132282 51128
rect 186314 51116 186320 51128
rect 132276 51088 186320 51116
rect 132276 51076 132282 51088
rect 186314 51076 186320 51088
rect 186372 51076 186378 51128
rect 132126 51008 132132 51060
rect 132184 51048 132190 51060
rect 137278 51048 137284 51060
rect 132184 51020 137284 51048
rect 132184 51008 132190 51020
rect 137278 51008 137284 51020
rect 137336 51008 137342 51060
rect 133506 49716 133512 49768
rect 133564 49756 133570 49768
rect 186314 49756 186320 49768
rect 133564 49728 186320 49756
rect 133564 49716 133570 49728
rect 186314 49716 186320 49728
rect 186372 49716 186378 49768
rect 131206 49648 131212 49700
rect 131264 49688 131270 49700
rect 148318 49688 148324 49700
rect 131264 49660 148324 49688
rect 131264 49648 131270 49660
rect 148318 49648 148324 49660
rect 148376 49648 148382 49700
rect 131298 49580 131304 49632
rect 131356 49620 131362 49632
rect 133230 49620 133236 49632
rect 131356 49592 133236 49620
rect 131356 49580 131362 49592
rect 133230 49580 133236 49592
rect 133288 49580 133294 49632
rect 131850 48288 131856 48340
rect 131908 48328 131914 48340
rect 186314 48328 186320 48340
rect 131908 48300 186320 48328
rect 131908 48288 131914 48300
rect 186314 48288 186320 48300
rect 186372 48288 186378 48340
rect 411254 48288 411260 48340
rect 411312 48328 411318 48340
rect 417510 48328 417516 48340
rect 411312 48300 417516 48328
rect 411312 48288 411318 48300
rect 417510 48288 417516 48300
rect 417568 48288 417574 48340
rect 131206 48220 131212 48272
rect 131264 48260 131270 48272
rect 187142 48260 187148 48272
rect 131264 48232 187148 48260
rect 131264 48220 131270 48232
rect 187142 48220 187148 48232
rect 187200 48220 187206 48272
rect 416314 48220 416320 48272
rect 416372 48260 416378 48272
rect 437474 48260 437480 48272
rect 416372 48232 437480 48260
rect 416372 48220 416378 48232
rect 437474 48220 437480 48232
rect 437532 48220 437538 48272
rect 132218 48152 132224 48204
rect 132276 48192 132282 48204
rect 146938 48192 146944 48204
rect 132276 48164 146944 48192
rect 132276 48152 132282 48164
rect 146938 48152 146944 48164
rect 146996 48152 147002 48204
rect 132494 46928 132500 46980
rect 132552 46968 132558 46980
rect 186314 46968 186320 46980
rect 132552 46940 186320 46968
rect 132552 46928 132558 46940
rect 186314 46928 186320 46940
rect 186372 46928 186378 46980
rect 131114 46860 131120 46912
rect 131172 46900 131178 46912
rect 144178 46900 144184 46912
rect 131172 46872 144184 46900
rect 131172 46860 131178 46872
rect 144178 46860 144184 46872
rect 144236 46860 144242 46912
rect 412266 46860 412272 46912
rect 412324 46900 412330 46912
rect 437474 46900 437480 46912
rect 412324 46872 437480 46900
rect 412324 46860 412330 46872
rect 437474 46860 437480 46872
rect 437532 46860 437538 46912
rect 131114 45500 131120 45552
rect 131172 45540 131178 45552
rect 133322 45540 133328 45552
rect 131172 45512 133328 45540
rect 131172 45500 131178 45512
rect 133322 45500 133328 45512
rect 133380 45500 133386 45552
rect 419166 45500 419172 45552
rect 419224 45540 419230 45552
rect 437474 45540 437480 45552
rect 419224 45512 437480 45540
rect 419224 45500 419230 45512
rect 437474 45500 437480 45512
rect 437532 45500 437538 45552
rect 131206 45432 131212 45484
rect 131264 45472 131270 45484
rect 187050 45472 187056 45484
rect 131264 45444 187056 45472
rect 131264 45432 131270 45444
rect 187050 45432 187056 45444
rect 187108 45432 187114 45484
rect 131206 44072 131212 44124
rect 131264 44112 131270 44124
rect 187234 44112 187240 44124
rect 131264 44084 187240 44112
rect 131264 44072 131270 44084
rect 187234 44072 187240 44084
rect 187292 44072 187298 44124
rect 416406 44072 416412 44124
rect 416464 44112 416470 44124
rect 437474 44112 437480 44124
rect 416464 44084 437480 44112
rect 416464 44072 416470 44084
rect 437474 44072 437480 44084
rect 437532 44072 437538 44124
rect 131666 42848 131672 42900
rect 131724 42888 131730 42900
rect 186406 42888 186412 42900
rect 131724 42860 186412 42888
rect 131724 42848 131730 42860
rect 186406 42848 186412 42860
rect 186464 42848 186470 42900
rect 131298 42780 131304 42832
rect 131356 42820 131362 42832
rect 186314 42820 186320 42832
rect 131356 42792 186320 42820
rect 131356 42780 131362 42792
rect 186314 42780 186320 42792
rect 186372 42780 186378 42832
rect 131114 42712 131120 42764
rect 131172 42752 131178 42764
rect 187326 42752 187332 42764
rect 131172 42724 187332 42752
rect 131172 42712 131178 42724
rect 187326 42712 187332 42724
rect 187384 42712 187390 42764
rect 411898 42712 411904 42764
rect 411956 42752 411962 42764
rect 437474 42752 437480 42764
rect 411956 42724 437480 42752
rect 411956 42712 411962 42724
rect 437474 42712 437480 42724
rect 437532 42712 437538 42764
rect 131206 42644 131212 42696
rect 131264 42684 131270 42696
rect 133414 42684 133420 42696
rect 131264 42656 133420 42684
rect 131264 42644 131270 42656
rect 133414 42644 133420 42656
rect 133472 42644 133478 42696
rect 411254 42644 411260 42696
rect 411312 42684 411318 42696
rect 414842 42684 414848 42696
rect 411312 42656 414848 42684
rect 411312 42644 411318 42656
rect 414842 42644 414848 42656
rect 414900 42644 414906 42696
rect 131114 41352 131120 41404
rect 131172 41392 131178 41404
rect 186958 41392 186964 41404
rect 131172 41364 186964 41392
rect 131172 41352 131178 41364
rect 186958 41352 186964 41364
rect 187016 41352 187022 41404
rect 417970 41352 417976 41404
rect 418028 41392 418034 41404
rect 437474 41392 437480 41404
rect 418028 41364 437480 41392
rect 418028 41352 418034 41364
rect 437474 41352 437480 41364
rect 437532 41352 437538 41404
rect 131206 41284 131212 41336
rect 131264 41324 131270 41336
rect 133506 41324 133512 41336
rect 131264 41296 133512 41324
rect 131264 41284 131270 41296
rect 133506 41284 133512 41296
rect 133564 41284 133570 41336
rect 411254 41012 411260 41064
rect 411312 41052 411318 41064
rect 414750 41052 414756 41064
rect 411312 41024 414756 41052
rect 411312 41012 411318 41024
rect 414750 41012 414756 41024
rect 414808 41012 414814 41064
rect 411898 40672 411904 40724
rect 411956 40712 411962 40724
rect 412174 40712 412180 40724
rect 411956 40684 412180 40712
rect 411956 40672 411962 40684
rect 412174 40672 412180 40684
rect 412232 40672 412238 40724
rect 411254 38836 411260 38888
rect 411312 38876 411318 38888
rect 414658 38876 414664 38888
rect 411312 38848 414664 38876
rect 411312 38836 411318 38848
rect 414658 38836 414664 38848
rect 414716 38836 414722 38888
rect 131206 38564 131212 38616
rect 131264 38604 131270 38616
rect 187142 38604 187148 38616
rect 131264 38576 187148 38604
rect 131264 38564 131270 38576
rect 187142 38564 187148 38576
rect 187200 38564 187206 38616
rect 416498 38564 416504 38616
rect 416556 38604 416562 38616
rect 437474 38604 437480 38616
rect 416556 38576 437480 38604
rect 416556 38564 416562 38576
rect 437474 38564 437480 38576
rect 437532 38564 437538 38616
rect 131114 38496 131120 38548
rect 131172 38536 131178 38548
rect 186590 38536 186596 38548
rect 131172 38508 186596 38536
rect 131172 38496 131178 38508
rect 186590 38496 186596 38508
rect 186648 38496 186654 38548
rect 132126 37340 132132 37392
rect 132184 37380 132190 37392
rect 186406 37380 186412 37392
rect 132184 37352 186412 37380
rect 132184 37340 132190 37352
rect 186406 37340 186412 37352
rect 186464 37340 186470 37392
rect 132034 37272 132040 37324
rect 132092 37312 132098 37324
rect 186314 37312 186320 37324
rect 132092 37284 186320 37312
rect 132092 37272 132098 37284
rect 186314 37272 186320 37284
rect 186372 37272 186378 37324
rect 131206 37204 131212 37256
rect 131264 37244 131270 37256
rect 186498 37244 186504 37256
rect 131264 37216 186504 37244
rect 131264 37204 131270 37216
rect 186498 37204 186504 37216
rect 186556 37204 186562 37256
rect 411990 37204 411996 37256
rect 412048 37244 412054 37256
rect 437474 37244 437480 37256
rect 412048 37216 437480 37244
rect 412048 37204 412054 37216
rect 437474 37204 437480 37216
rect 437532 37204 437538 37256
rect 411254 37136 411260 37188
rect 411312 37176 411318 37188
rect 438210 37176 438216 37188
rect 411312 37148 438216 37176
rect 411312 37136 411318 37148
rect 438210 37136 438216 37148
rect 438268 37136 438274 37188
rect 132218 35912 132224 35964
rect 132276 35952 132282 35964
rect 186314 35952 186320 35964
rect 132276 35924 186320 35952
rect 132276 35912 132282 35924
rect 186314 35912 186320 35924
rect 186372 35912 186378 35964
rect 131206 35844 131212 35896
rect 131264 35884 131270 35896
rect 187234 35884 187240 35896
rect 131264 35856 187240 35884
rect 131264 35844 131270 35856
rect 187234 35844 187240 35856
rect 187292 35844 187298 35896
rect 416038 35844 416044 35896
rect 416096 35884 416102 35896
rect 437474 35884 437480 35896
rect 416096 35856 437480 35884
rect 416096 35844 416102 35856
rect 437474 35844 437480 35856
rect 437532 35844 437538 35896
rect 131114 35776 131120 35828
rect 131172 35816 131178 35828
rect 186958 35816 186964 35828
rect 131172 35788 186964 35816
rect 131172 35776 131178 35788
rect 186958 35776 186964 35788
rect 187016 35776 187022 35828
rect 411254 35776 411260 35828
rect 411312 35816 411318 35828
rect 418890 35816 418896 35828
rect 411312 35788 418896 35816
rect 411312 35776 411318 35788
rect 418890 35776 418896 35788
rect 418948 35776 418954 35828
rect 415118 34416 415124 34468
rect 415176 34456 415182 34468
rect 437474 34456 437480 34468
rect 415176 34428 437480 34456
rect 415176 34416 415182 34428
rect 437474 34416 437480 34428
rect 437532 34416 437538 34468
rect 131114 33124 131120 33176
rect 131172 33164 131178 33176
rect 186314 33164 186320 33176
rect 131172 33136 186320 33164
rect 131172 33124 131178 33136
rect 186314 33124 186320 33136
rect 186372 33124 186378 33176
rect 131206 33056 131212 33108
rect 131264 33096 131270 33108
rect 186406 33096 186412 33108
rect 131264 33068 186412 33096
rect 131264 33056 131270 33068
rect 186406 33056 186412 33068
rect 186464 33056 186470 33108
rect 411254 33056 411260 33108
rect 411312 33096 411318 33108
rect 438118 33096 438124 33108
rect 411312 33068 438124 33096
rect 411312 33056 411318 33068
rect 438118 33056 438124 33068
rect 438176 33056 438182 33108
rect 412082 32988 412088 33040
rect 412140 33028 412146 33040
rect 437474 33028 437480 33040
rect 412140 33000 437480 33028
rect 412140 32988 412146 33000
rect 437474 32988 437480 33000
rect 437532 32988 437538 33040
rect 131298 31832 131304 31884
rect 131356 31872 131362 31884
rect 186314 31872 186320 31884
rect 131356 31844 186320 31872
rect 131356 31832 131362 31844
rect 186314 31832 186320 31844
rect 186372 31832 186378 31884
rect 131206 31764 131212 31816
rect 131264 31804 131270 31816
rect 186406 31804 186412 31816
rect 131264 31776 186412 31804
rect 131264 31764 131270 31776
rect 186406 31764 186412 31776
rect 186464 31764 186470 31816
rect 412266 31696 412272 31748
rect 412324 31736 412330 31748
rect 542630 31736 542636 31748
rect 412324 31708 542636 31736
rect 412324 31696 412330 31708
rect 542630 31696 542636 31708
rect 542688 31696 542694 31748
rect 412542 31628 412548 31680
rect 412600 31668 412606 31680
rect 542538 31668 542544 31680
rect 412600 31640 542544 31668
rect 412600 31628 412606 31640
rect 542538 31628 542544 31640
rect 542596 31628 542602 31680
rect 412358 31560 412364 31612
rect 412416 31600 412422 31612
rect 437474 31600 437480 31612
rect 412416 31572 437480 31600
rect 412416 31560 412422 31572
rect 437474 31560 437480 31572
rect 437532 31560 437538 31612
rect 131114 31016 131120 31068
rect 131172 31056 131178 31068
rect 186314 31056 186320 31068
rect 131172 31028 186320 31056
rect 131172 31016 131178 31028
rect 186314 31016 186320 31028
rect 186372 31016 186378 31068
rect 186682 30268 186688 30320
rect 186740 30308 186746 30320
rect 580166 30308 580172 30320
rect 186740 30280 580172 30308
rect 186740 30268 186746 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 411254 30200 411260 30252
rect 411312 30240 411318 30252
rect 542722 30240 542728 30252
rect 411312 30212 542728 30240
rect 411312 30200 411318 30212
rect 542722 30200 542728 30212
rect 542780 30200 542786 30252
rect 411898 30132 411904 30184
rect 411956 30172 411962 30184
rect 542354 30172 542360 30184
rect 411956 30144 542360 30172
rect 411956 30132 411962 30144
rect 542354 30132 542360 30144
rect 542412 30132 542418 30184
rect 412450 30064 412456 30116
rect 412508 30104 412514 30116
rect 542446 30104 542452 30116
rect 412508 30076 542452 30104
rect 412508 30064 412514 30076
rect 542446 30064 542452 30076
rect 542504 30064 542510 30116
rect 188430 29452 188436 29504
rect 188488 29492 188494 29504
rect 258902 29492 258908 29504
rect 188488 29464 258908 29492
rect 188488 29452 188494 29464
rect 258902 29452 258908 29464
rect 258960 29452 258966 29504
rect 188522 29384 188528 29436
rect 188580 29424 188586 29436
rect 299566 29424 299572 29436
rect 188580 29396 299572 29424
rect 188580 29384 188586 29396
rect 299566 29384 299572 29396
rect 299624 29384 299630 29436
rect 130470 29316 130476 29368
rect 130528 29356 130534 29368
rect 242986 29356 242992 29368
rect 130528 29328 242992 29356
rect 130528 29316 130534 29328
rect 242986 29316 242992 29328
rect 243044 29316 243050 29368
rect 417510 29316 417516 29368
rect 417568 29356 417574 29368
rect 468754 29356 468760 29368
rect 417568 29328 468760 29356
rect 417568 29316 417574 29328
rect 468754 29316 468760 29328
rect 468812 29316 468818 29368
rect 201494 29248 201500 29300
rect 201552 29288 201558 29300
rect 202506 29288 202512 29300
rect 201552 29260 202512 29288
rect 201552 29248 201558 29260
rect 202506 29248 202512 29260
rect 202564 29288 202570 29300
rect 410610 29288 410616 29300
rect 202564 29260 410616 29288
rect 202564 29248 202570 29260
rect 410610 29248 410616 29260
rect 410668 29248 410674 29300
rect 413462 29248 413468 29300
rect 413520 29288 413526 29300
rect 485774 29288 485780 29300
rect 413520 29260 485780 29288
rect 413520 29248 413526 29260
rect 485774 29248 485780 29260
rect 485832 29248 485838 29300
rect 193214 29180 193220 29232
rect 193272 29220 193278 29232
rect 194410 29220 194416 29232
rect 193272 29192 194416 29220
rect 193272 29180 193278 29192
rect 194410 29180 194416 29192
rect 194468 29220 194474 29232
rect 410518 29220 410524 29232
rect 194468 29192 410524 29220
rect 194468 29180 194474 29192
rect 410518 29180 410524 29192
rect 410576 29180 410582 29232
rect 452562 29180 452568 29232
rect 452620 29220 452626 29232
rect 580350 29220 580356 29232
rect 452620 29192 580356 29220
rect 452620 29180 452626 29192
rect 580350 29180 580356 29192
rect 580408 29180 580414 29232
rect 130378 29112 130384 29164
rect 130436 29152 130442 29164
rect 364702 29152 364708 29164
rect 130436 29124 364708 29152
rect 130436 29112 130442 29124
rect 364702 29112 364708 29124
rect 364760 29112 364766 29164
rect 444282 29112 444288 29164
rect 444340 29152 444346 29164
rect 580258 29152 580264 29164
rect 444340 29124 580264 29152
rect 444340 29112 444346 29124
rect 580258 29112 580264 29124
rect 580316 29112 580322 29164
rect 226978 29044 226984 29096
rect 227036 29084 227042 29096
rect 580442 29084 580448 29096
rect 227036 29056 580448 29084
rect 227036 29044 227042 29056
rect 580442 29044 580448 29056
rect 580500 29044 580506 29096
rect 210602 28976 210608 29028
rect 210660 29016 210666 29028
rect 580534 29016 580540 29028
rect 210660 28988 580540 29016
rect 210660 28976 210666 28988
rect 580534 28976 580540 28988
rect 580592 28976 580598 29028
rect 130562 28908 130568 28960
rect 130620 28948 130626 28960
rect 381078 28948 381084 28960
rect 130620 28920 381084 28948
rect 130620 28908 130626 28920
rect 381078 28908 381084 28920
rect 381136 28908 381142 28960
rect 413370 28908 413376 28960
rect 413428 28948 413434 28960
rect 535454 28948 535460 28960
rect 413428 28920 535460 28948
rect 413428 28908 413434 28920
rect 535454 28908 535460 28920
rect 535512 28908 535518 28960
rect 130654 28840 130660 28892
rect 130712 28880 130718 28892
rect 372982 28880 372988 28892
rect 130712 28852 372988 28880
rect 130712 28840 130718 28852
rect 372982 28840 372988 28852
rect 373040 28840 373046 28892
rect 418982 28840 418988 28892
rect 419040 28880 419046 28892
rect 518986 28880 518992 28892
rect 419040 28852 518992 28880
rect 419040 28840 419046 28852
rect 518986 28840 518992 28852
rect 519044 28840 519050 28892
rect 188706 28772 188712 28824
rect 188764 28812 188770 28824
rect 389174 28812 389180 28824
rect 188764 28784 389180 28812
rect 188764 28772 188770 28784
rect 389174 28772 389180 28784
rect 389232 28772 389238 28824
rect 439498 28772 439504 28824
rect 439556 28812 439562 28824
rect 527174 28812 527180 28824
rect 439556 28784 527180 28812
rect 439556 28772 439562 28784
rect 527174 28772 527180 28784
rect 527232 28772 527238 28824
rect 188890 28704 188896 28756
rect 188948 28744 188954 28756
rect 356606 28744 356612 28756
rect 188948 28716 356612 28744
rect 188948 28704 188954 28716
rect 356606 28704 356612 28716
rect 356664 28704 356670 28756
rect 417418 28704 417424 28756
rect 417476 28744 417482 28756
rect 502334 28744 502340 28756
rect 417476 28716 502340 28744
rect 417476 28704 417482 28716
rect 502334 28704 502340 28716
rect 502392 28704 502398 28756
rect 188982 28636 188988 28688
rect 189040 28676 189046 28688
rect 348510 28676 348516 28688
rect 189040 28648 348516 28676
rect 189040 28636 189046 28648
rect 348510 28636 348516 28648
rect 348568 28636 348574 28688
rect 436738 28636 436744 28688
rect 436796 28676 436802 28688
rect 510614 28676 510620 28688
rect 436796 28648 510620 28676
rect 436796 28636 436802 28648
rect 510614 28636 510620 28648
rect 510672 28636 510678 28688
rect 182818 28568 182824 28620
rect 182876 28608 182882 28620
rect 340414 28608 340420 28620
rect 182876 28580 340420 28608
rect 182876 28568 182882 28580
rect 340414 28568 340420 28580
rect 340472 28568 340478 28620
rect 413278 28568 413284 28620
rect 413336 28608 413342 28620
rect 477494 28608 477500 28620
rect 413336 28580 477500 28608
rect 413336 28568 413342 28580
rect 477494 28568 477500 28580
rect 477552 28568 477558 28620
rect 188154 28500 188160 28552
rect 188212 28540 188218 28552
rect 332134 28540 332140 28552
rect 188212 28512 332140 28540
rect 188212 28500 188218 28512
rect 332134 28500 332140 28512
rect 332192 28500 332198 28552
rect 439590 28500 439596 28552
rect 439648 28540 439654 28552
rect 494146 28540 494152 28552
rect 439648 28512 494152 28540
rect 439648 28500 439654 28512
rect 494146 28500 494152 28512
rect 494204 28500 494210 28552
rect 188246 28432 188252 28484
rect 188304 28472 188310 28484
rect 324406 28472 324412 28484
rect 188304 28444 324412 28472
rect 188304 28432 188310 28444
rect 324406 28432 324412 28444
rect 324464 28432 324470 28484
rect 188798 28364 188804 28416
rect 188856 28404 188862 28416
rect 316126 28404 316132 28416
rect 188856 28376 316132 28404
rect 188856 28364 188862 28376
rect 316126 28364 316132 28376
rect 316184 28364 316190 28416
rect 189810 28296 189816 28348
rect 189868 28336 189874 28348
rect 307754 28336 307760 28348
rect 189868 28308 307760 28336
rect 189868 28296 189874 28308
rect 307754 28296 307760 28308
rect 307812 28296 307818 28348
rect 188614 28228 188620 28280
rect 188672 28268 188678 28280
rect 283374 28268 283380 28280
rect 188672 28240 283380 28268
rect 188672 28228 188678 28240
rect 283374 28228 283380 28240
rect 283432 28228 283438 28280
rect 189902 28160 189908 28212
rect 189960 28200 189966 28212
rect 275094 28200 275100 28212
rect 189960 28172 275100 28200
rect 189960 28160 189966 28172
rect 275094 28160 275100 28172
rect 275152 28160 275158 28212
rect 189718 28092 189724 28144
rect 189776 28132 189782 28144
rect 266998 28132 267004 28144
rect 189776 28104 267004 28132
rect 189776 28092 189782 28104
rect 266998 28092 267004 28104
rect 267056 28092 267062 28144
rect 188338 28024 188344 28076
rect 188396 28064 188402 28076
rect 234614 28064 234620 28076
rect 188396 28036 234620 28064
rect 188396 28024 188402 28036
rect 234614 28024 234620 28036
rect 234672 28024 234678 28076
rect 79962 27548 79968 27600
rect 80020 27588 80026 27600
rect 460474 27588 460480 27600
rect 80020 27560 460480 27588
rect 80020 27548 80026 27560
rect 460474 27548 460480 27560
rect 460532 27548 460538 27600
rect 418798 20612 418804 20664
rect 418856 20652 418862 20664
rect 579982 20652 579988 20664
rect 418856 20624 579988 20652
rect 418856 20612 418862 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 218054 6808 218060 6860
rect 218112 6848 218118 6860
rect 580166 6848 580172 6860
rect 218112 6820 580172 6848
rect 218112 6808 218118 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 2682 4088 2688 4140
rect 2740 4128 2746 4140
rect 201494 4128 201500 4140
rect 2740 4100 201500 4128
rect 2740 4088 2746 4100
rect 201494 4088 201500 4100
rect 201552 4088 201558 4140
rect 1302 4020 1308 4072
rect 1360 4060 1366 4072
rect 193214 4060 193220 4072
rect 1360 4032 193220 4060
rect 1360 4020 1366 4032
rect 193214 4020 193220 4032
rect 193272 4020 193278 4072
rect 1670 3680 1676 3732
rect 1728 3720 1734 3732
rect 2682 3720 2688 3732
rect 1728 3692 2688 3720
rect 1728 3680 1734 3692
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 566 3612 572 3664
rect 624 3652 630 3664
rect 1302 3652 1308 3664
rect 624 3624 1308 3652
rect 624 3612 630 3624
rect 1302 3612 1308 3624
rect 1360 3612 1366 3664
<< via1 >>
rect 204260 325660 204312 325712
rect 207020 325660 207072 325712
rect 193220 306348 193272 306400
rect 207020 306348 207072 306400
rect 190460 304988 190512 305040
rect 207020 304988 207072 305040
rect 55220 298120 55272 298172
rect 55864 298120 55916 298172
rect 215852 298120 215904 298172
rect 95148 297508 95200 297560
rect 130384 297508 130436 297560
rect 71504 297440 71556 297492
rect 130476 297440 130528 297492
rect 81808 297372 81860 297424
rect 188528 297372 188580 297424
rect 76840 297304 76892 297356
rect 188436 297304 188488 297356
rect 65708 297236 65760 297288
rect 188344 297236 188396 297288
rect 67824 297168 67876 297220
rect 227720 297168 227772 297220
rect 70216 297100 70268 297152
rect 229100 297100 229152 297152
rect 229468 297100 229520 297152
rect 69940 297032 69992 297084
rect 229192 297032 229244 297084
rect 79784 296964 79836 297016
rect 352564 296964 352616 297016
rect 106740 296896 106792 296948
rect 409144 296896 409196 296948
rect 103244 296828 103296 296880
rect 409052 296828 409104 296880
rect 96712 296760 96764 296812
rect 408960 296760 409012 296812
rect 93308 296692 93360 296744
rect 408868 296692 408920 296744
rect 267464 263236 267516 263288
rect 371332 263236 371384 263288
rect 110328 263168 110380 263220
rect 411628 263168 411680 263220
rect 104716 263100 104768 263152
rect 410432 263100 410484 263152
rect 99196 263032 99248 263084
rect 411536 263032 411588 263084
rect 86684 262964 86736 263016
rect 409972 262964 410024 263016
rect 81256 262896 81308 262948
rect 410064 262896 410116 262948
rect 75828 262828 75880 262880
rect 411720 262828 411772 262880
rect 259184 261876 259236 261928
rect 338120 261876 338172 261928
rect 263416 261808 263468 261860
rect 352104 261808 352156 261860
rect 264796 261740 264848 261792
rect 356704 261740 356756 261792
rect 266176 261672 266228 261724
rect 361580 261672 361632 261724
rect 267556 261604 267608 261656
rect 366088 261604 366140 261656
rect 104808 261536 104860 261588
rect 406016 261536 406068 261588
rect 81348 261468 81400 261520
rect 385040 261468 385092 261520
rect 253756 260584 253808 260636
rect 314752 260584 314804 260636
rect 255136 260516 255188 260568
rect 319352 260516 319404 260568
rect 256516 260448 256568 260500
rect 324320 260448 324372 260500
rect 257804 260380 257856 260432
rect 328736 260380 328788 260432
rect 259276 260312 259328 260364
rect 333336 260312 333388 260364
rect 260656 260244 260708 260296
rect 342720 260244 342772 260296
rect 79876 260176 79928 260228
rect 378140 260176 378192 260228
rect 100576 260108 100628 260160
rect 401600 260108 401652 260160
rect 246764 259020 246816 259072
rect 286600 259020 286652 259072
rect 248236 258952 248288 259004
rect 291200 258952 291252 259004
rect 249616 258884 249668 258936
rect 295984 258884 296036 258936
rect 250996 258816 251048 258868
rect 300860 258816 300912 258868
rect 252284 258748 252336 258800
rect 305368 258748 305420 258800
rect 262036 258680 262088 258732
rect 347780 258680 347832 258732
rect 245568 257796 245620 257848
rect 282092 257796 282144 257848
rect 260748 257728 260800 257780
rect 307760 257728 307812 257780
rect 262128 257660 262180 257712
rect 312452 257660 312504 257712
rect 263508 257592 263560 257644
rect 317512 257592 317564 257644
rect 266268 257524 266320 257576
rect 326436 257524 326488 257576
rect 273076 257456 273128 257508
rect 354772 257456 354824 257508
rect 90916 257388 90968 257440
rect 410340 257388 410392 257440
rect 78496 257320 78548 257372
rect 409880 257320 409932 257372
rect 242808 256504 242860 256556
rect 268016 256504 268068 256556
rect 255228 256436 255280 256488
rect 284300 256436 284352 256488
rect 219256 256368 219308 256420
rect 229192 256368 229244 256420
rect 256608 256368 256660 256420
rect 289084 256368 289136 256420
rect 210056 256300 210108 256352
rect 227720 256300 227772 256352
rect 257896 256300 257948 256352
rect 293960 256300 294012 256352
rect 212448 256232 212500 256284
rect 231860 256232 231912 256284
rect 257988 256232 258040 256284
rect 298468 256232 298520 256284
rect 201408 256164 201460 256216
rect 226340 256164 226392 256216
rect 259368 256164 259420 256216
rect 303068 256164 303120 256216
rect 93676 256096 93728 256148
rect 250352 256096 250404 256148
rect 277308 256096 277360 256148
rect 368572 256096 368624 256148
rect 49608 256028 49660 256080
rect 387340 256028 387392 256080
rect 47952 255960 48004 256012
rect 410248 255960 410300 256012
rect 217048 255008 217100 255060
rect 240140 255008 240192 255060
rect 252468 255008 252520 255060
rect 274916 255008 274968 255060
rect 202696 254940 202748 254992
rect 230480 254940 230532 254992
rect 253848 254940 253900 254992
rect 279700 254940 279752 254992
rect 209596 254872 209648 254924
rect 240140 254872 240192 254924
rect 244096 254872 244148 254924
rect 277492 254872 277544 254924
rect 207848 254804 207900 254856
rect 238760 254804 238812 254856
rect 252376 254804 252428 254856
rect 310060 254804 310112 254856
rect 209688 254736 209740 254788
rect 247040 254736 247092 254788
rect 251088 254736 251140 254788
rect 270500 254736 270552 254788
rect 273168 254736 273220 254788
rect 349804 254736 349856 254788
rect 47676 254668 47728 254720
rect 373356 254668 373408 254720
rect 47768 254600 47820 254652
rect 382556 254600 382608 254652
rect 47860 254532 47912 254584
rect 410156 254532 410208 254584
rect 228732 253852 228784 253904
rect 229100 253852 229152 253904
rect 246948 253852 247000 253904
rect 249156 253852 249208 253904
rect 242808 253784 242860 253836
rect 244280 253784 244332 253836
rect 264888 253580 264940 253632
rect 321836 253580 321888 253632
rect 208032 253512 208084 253564
rect 214196 253512 214248 253564
rect 221832 253512 221884 253564
rect 233240 253512 233292 253564
rect 237196 253512 237248 253564
rect 244556 253512 244608 253564
rect 246856 253512 246908 253564
rect 256332 253512 256384 253564
rect 267648 253512 267700 253564
rect 331220 253512 331272 253564
rect 208124 253444 208176 253496
rect 223580 253444 223632 253496
rect 226248 253444 226300 253496
rect 241520 253444 241572 253496
rect 248328 253444 248380 253496
rect 260932 253444 260984 253496
rect 269028 253444 269080 253496
rect 335820 253444 335872 253496
rect 208216 253376 208268 253428
rect 232780 253376 232832 253428
rect 235816 253376 235868 253428
rect 242900 253376 242952 253428
rect 249708 253376 249760 253428
rect 265532 253376 265584 253428
rect 270408 253376 270460 253428
rect 340420 253376 340472 253428
rect 195796 253308 195848 253360
rect 224960 253308 225012 253360
rect 240048 253308 240100 253360
rect 258540 253308 258592 253360
rect 271788 253308 271840 253360
rect 345204 253308 345256 253360
rect 198464 253240 198516 253292
rect 237380 253240 237432 253292
rect 244188 253240 244240 253292
rect 272708 253240 272760 253292
rect 274548 253240 274600 253292
rect 359188 253240 359240 253292
rect 77116 253172 77168 253224
rect 147680 253172 147732 253224
rect 208308 253172 208360 253224
rect 253940 253172 253992 253224
rect 275928 253172 275980 253224
rect 363972 253172 364024 253224
rect 231216 253104 231268 253156
rect 234620 253104 234672 253156
rect 67548 252492 67600 252544
rect 200488 252492 200540 252544
rect 201408 252492 201460 252544
rect 238668 252356 238720 252408
rect 251548 252356 251600 252408
rect 241428 252288 241480 252340
rect 263692 252288 263744 252340
rect 352564 252288 352616 252340
rect 394332 252288 394384 252340
rect 250352 252220 250404 252272
rect 403716 252220 403768 252272
rect 147680 252152 147732 252204
rect 391940 252152 391992 252204
rect 111708 252084 111760 252136
rect 408592 252084 408644 252136
rect 84016 252016 84068 252068
rect 389732 252016 389784 252068
rect 91008 251948 91060 252000
rect 398932 251948 398984 252000
rect 88156 251880 88208 251932
rect 396724 251880 396776 251932
rect 49516 251812 49568 251864
rect 375564 251812 375616 251864
rect 117228 250792 117280 250844
rect 408500 250792 408552 250844
rect 114468 250724 114520 250776
rect 410524 250724 410576 250776
rect 115848 250656 115900 250708
rect 411260 250656 411312 250708
rect 107476 250588 107528 250640
rect 411444 250588 411496 250640
rect 73068 250520 73120 250572
rect 411812 250520 411864 250572
rect 48044 250452 48096 250504
rect 411352 250452 411404 250504
rect 187240 249772 187292 249824
rect 580356 249772 580408 249824
rect 106096 249704 106148 249756
rect 187516 249704 187568 249756
rect 108856 249636 108908 249688
rect 187608 249636 187660 249688
rect 187424 248412 187476 248464
rect 580264 248412 580316 248464
rect 112996 248344 113048 248396
rect 187608 248344 187660 248396
rect 113088 246984 113140 247036
rect 187332 246984 187384 247036
rect 101864 245556 101916 245608
rect 187608 245556 187660 245608
rect 101956 244196 102008 244248
rect 186320 244196 186372 244248
rect 411260 243516 411312 243568
rect 411444 243516 411496 243568
rect 411444 243380 411496 243432
rect 411812 243380 411864 243432
rect 102048 242836 102100 242888
rect 186412 242836 186464 242888
rect 106188 242768 106240 242820
rect 186320 242768 186372 242820
rect 93584 241408 93636 241460
rect 186320 241408 186372 241460
rect 99288 240048 99340 240100
rect 186320 240048 186372 240100
rect 89536 238688 89588 238740
rect 186320 238688 186372 238740
rect 86776 237328 86828 237380
rect 186412 237328 186464 237380
rect 96436 237260 96488 237312
rect 186320 237260 186372 237312
rect 95056 235900 95108 235952
rect 186320 235900 186372 235952
rect 89628 234540 89680 234592
rect 186320 234540 186372 234592
rect 78588 233180 78640 233232
rect 186320 233180 186372 233232
rect 463700 231820 463752 231872
rect 579620 231820 579672 231872
rect 48136 231752 48188 231804
rect 186320 231752 186372 231804
rect 82636 230392 82688 230444
rect 186320 230392 186372 230444
rect 74448 229032 74500 229084
rect 186320 229032 186372 229084
rect 169024 222164 169076 222216
rect 186320 222164 186372 222216
rect 131856 220804 131908 220856
rect 186320 220804 186372 220856
rect 159364 219444 159416 219496
rect 186320 219444 186372 219496
rect 135996 218016 136048 218068
rect 186320 218016 186372 218068
rect 543004 218016 543056 218068
rect 580172 218016 580224 218068
rect 142804 216724 142856 216776
rect 186412 216724 186464 216776
rect 135904 216656 135956 216708
rect 186320 216656 186372 216708
rect 157984 215296 158036 215348
rect 186320 215296 186372 215348
rect 134524 213936 134576 213988
rect 186320 213936 186372 213988
rect 141424 212508 141476 212560
rect 186320 212508 186372 212560
rect 156604 211148 156656 211200
rect 186320 211148 186372 211200
rect 136088 209788 136140 209840
rect 186320 209788 186372 209840
rect 411260 209788 411312 209840
rect 418804 209788 418856 209840
rect 141516 208360 141568 208412
rect 186320 208360 186372 208412
rect 133236 207000 133288 207052
rect 186320 207000 186372 207052
rect 411260 207000 411312 207052
rect 414664 207000 414716 207052
rect 155224 205640 155276 205692
rect 186320 205640 186372 205692
rect 411260 205640 411312 205692
rect 544384 205640 544436 205692
rect 142896 204280 142948 204332
rect 186320 204280 186372 204332
rect 134616 202852 134668 202904
rect 186320 202852 186372 202904
rect 411260 202852 411312 202904
rect 540244 202852 540296 202904
rect 152464 201492 152516 201544
rect 186320 201492 186372 201544
rect 134708 200132 134760 200184
rect 186320 200132 186372 200184
rect 151084 198772 151136 198824
rect 186412 198772 186464 198824
rect 134800 198704 134852 198756
rect 186320 198704 186372 198756
rect 148324 197344 148376 197396
rect 186320 197344 186372 197396
rect 411260 197344 411312 197396
rect 421564 197344 421616 197396
rect 134892 195984 134944 196036
rect 186320 195984 186372 196036
rect 411260 195984 411312 196036
rect 416044 195984 416096 196036
rect 145564 194556 145616 194608
rect 186320 194556 186372 194608
rect 134984 193196 135036 193248
rect 186320 193196 186372 193248
rect 146944 191904 146996 191956
rect 186412 191904 186464 191956
rect 133328 191836 133380 191888
rect 186320 191836 186372 191888
rect 411260 191836 411312 191888
rect 436744 191836 436796 191888
rect 543188 191836 543240 191888
rect 580172 191836 580224 191888
rect 147036 190476 147088 190528
rect 186320 190476 186372 190528
rect 145656 189048 145708 189100
rect 186320 189048 186372 189100
rect 411260 189048 411312 189100
rect 421656 189048 421708 189100
rect 140136 187688 140188 187740
rect 186320 187688 186372 187740
rect 411260 187688 411312 187740
rect 435364 187688 435416 187740
rect 140044 186396 140096 186448
rect 186320 186396 186372 186448
rect 133420 186328 133472 186380
rect 186412 186328 186464 186380
rect 411260 184900 411312 184952
rect 416136 184900 416188 184952
rect 137284 183540 137336 183592
rect 186320 183540 186372 183592
rect 411260 183540 411312 183592
rect 432604 183540 432656 183592
rect 145748 182180 145800 182232
rect 186320 182180 186372 182232
rect 411260 182180 411312 182232
rect 431224 182180 431276 182232
rect 140228 180820 140280 180872
rect 186320 180820 186372 180872
rect 140320 179460 140372 179512
rect 186320 179460 186372 179512
rect 133604 179392 133656 179444
rect 186412 179392 186464 179444
rect 411260 179392 411312 179444
rect 429844 179392 429896 179444
rect 133512 178032 133564 178084
rect 186320 178032 186372 178084
rect 411260 178032 411312 178084
rect 428464 178032 428516 178084
rect 543096 178032 543148 178084
rect 580172 178032 580224 178084
rect 138664 176672 138716 176724
rect 186320 176672 186372 176724
rect 133696 175244 133748 175296
rect 186320 175244 186372 175296
rect 411260 175244 411312 175296
rect 425704 175244 425756 175296
rect 137376 173884 137428 173936
rect 186320 173884 186372 173936
rect 411260 173884 411312 173936
rect 424324 173884 424376 173936
rect 138756 172524 138808 172576
rect 186320 172524 186372 172576
rect 411260 172524 411312 172576
rect 421748 172524 421800 172576
rect 145840 171096 145892 171148
rect 186320 171096 186372 171148
rect 166264 169736 166316 169788
rect 186320 169736 186372 169788
rect 411260 169736 411312 169788
rect 418988 169736 419040 169788
rect 136180 168376 136232 168428
rect 186320 168376 186372 168428
rect 411260 168376 411312 168428
rect 420276 168376 420328 168428
rect 138848 167084 138900 167136
rect 186320 167084 186372 167136
rect 131948 167016 132000 167068
rect 186412 167016 186464 167068
rect 164884 165588 164936 165640
rect 186320 165588 186372 165640
rect 411260 165588 411312 165640
rect 417424 165588 417476 165640
rect 138940 164228 138992 164280
rect 186320 164228 186372 164280
rect 411260 164228 411312 164280
rect 420184 164228 420236 164280
rect 132040 162868 132092 162920
rect 186320 162868 186372 162920
rect 162124 161508 162176 161560
rect 186320 161508 186372 161560
rect 135076 161440 135128 161492
rect 186412 161440 186464 161492
rect 411260 161440 411312 161492
rect 417608 161440 417660 161492
rect 136272 160080 136324 160132
rect 186320 160080 186372 160132
rect 411260 160080 411312 160132
rect 420368 160080 420420 160132
rect 132132 158720 132184 158772
rect 186320 158720 186372 158772
rect 411260 158720 411312 158772
rect 417516 158720 417568 158772
rect 139032 157360 139084 157412
rect 186320 157360 186372 157412
rect 160744 155932 160796 155984
rect 186320 155932 186372 155984
rect 411260 155932 411312 155984
rect 419080 155932 419132 155984
rect 137468 154640 137520 154692
rect 186320 154640 186372 154692
rect 133788 154572 133840 154624
rect 186412 154572 186464 154624
rect 411260 154572 411312 154624
rect 417700 154572 417752 154624
rect 145932 153212 145984 153264
rect 186320 153212 186372 153264
rect 147128 151784 147180 151836
rect 186320 151784 186372 151836
rect 411260 151784 411312 151836
rect 414940 151784 414992 151836
rect 146024 150424 146076 150476
rect 186320 150424 186372 150476
rect 411260 150424 411312 150476
rect 417792 150424 417844 150476
rect 144184 149132 144236 149184
rect 186320 149132 186372 149184
rect 137560 149064 137612 149116
rect 186412 149064 186464 149116
rect 132224 147636 132276 147688
rect 186320 147636 186372 147688
rect 411260 147636 411312 147688
rect 415032 147636 415084 147688
rect 144276 146276 144328 146328
rect 186320 146276 186372 146328
rect 411260 146276 411312 146328
rect 421840 146276 421892 146328
rect 143080 144916 143132 144968
rect 186320 144916 186372 144968
rect 411260 144916 411312 144968
rect 417884 144916 417936 144968
rect 141608 143556 141660 143608
rect 186320 143556 186372 143608
rect 144368 142196 144420 142248
rect 186412 142196 186464 142248
rect 142988 142128 143040 142180
rect 186320 142128 186372 142180
rect 411260 142128 411312 142180
rect 429936 142128 429988 142180
rect 411260 140768 411312 140820
rect 421932 140768 421984 140820
rect 137652 139408 137704 139460
rect 186320 139408 186372 139460
rect 414664 139340 414716 139392
rect 580172 139340 580224 139392
rect 143172 137980 143224 138032
rect 186320 137980 186372 138032
rect 411260 137980 411312 138032
rect 431316 137980 431368 138032
rect 141700 136620 141752 136672
rect 186320 136620 186372 136672
rect 411260 136620 411312 136672
rect 422024 136620 422076 136672
rect 143264 135328 143316 135380
rect 186320 135328 186372 135380
rect 137744 135260 137796 135312
rect 186412 135260 186464 135312
rect 140412 133900 140464 133952
rect 186320 133900 186372 133952
rect 411260 133900 411312 133952
rect 432696 133900 432748 133952
rect 137836 132472 137888 132524
rect 186320 132472 186372 132524
rect 411260 132472 411312 132524
rect 420460 132472 420512 132524
rect 103336 132268 103388 132320
rect 133144 132268 133196 132320
rect 100668 132200 100720 132252
rect 131672 132200 131724 132252
rect 97724 132132 97776 132184
rect 130568 132132 130620 132184
rect 108948 132064 109000 132116
rect 188712 132064 188764 132116
rect 97816 131996 97868 132048
rect 188988 131996 189040 132048
rect 88248 131928 88300 131980
rect 182824 131928 182876 131980
rect 92388 131860 92440 131912
rect 188804 131860 188856 131912
rect 92296 131792 92348 131844
rect 188896 131792 188948 131844
rect 48228 131724 48280 131776
rect 188620 131724 188672 131776
rect 419356 131452 419408 131504
rect 534632 131452 534684 131504
rect 410524 131384 410576 131436
rect 444656 131384 444708 131436
rect 414664 131316 414716 131368
rect 484584 131316 484636 131368
rect 414756 131248 414808 131300
rect 494612 131248 494664 131300
rect 1308 131180 1360 131232
rect 55128 131180 55180 131232
rect 414848 131180 414900 131232
rect 504640 131180 504692 131232
rect 2688 131112 2740 131164
rect 104900 131112 104952 131164
rect 141884 131112 141936 131164
rect 186320 131112 186372 131164
rect 96528 130704 96580 130756
rect 130660 130704 130712 130756
rect 85488 130636 85540 130688
rect 188252 130636 188304 130688
rect 85396 130568 85448 130620
rect 188160 130568 188212 130620
rect 86868 130500 86920 130552
rect 189816 130500 189868 130552
rect 85304 130432 85356 130484
rect 189724 130432 189776 130484
rect 84108 130364 84160 130416
rect 189816 130364 189868 130416
rect 434628 130364 434680 130416
rect 454592 130364 454644 130416
rect 418896 130024 418948 130076
rect 474740 130024 474792 130076
rect 413284 129956 413336 130008
rect 514760 129956 514812 130008
rect 413468 129888 413520 129940
rect 524604 129888 524656 129940
rect 415216 129820 415268 129872
rect 539324 129820 539376 129872
rect 144460 129752 144512 129804
rect 186320 129752 186372 129804
rect 413376 129752 413428 129804
rect 542452 129752 542504 129804
rect 131120 129684 131172 129736
rect 169024 129684 169076 129736
rect 131212 129616 131264 129668
rect 159364 129616 159416 129668
rect 411260 128460 411312 128512
rect 420552 128460 420604 128512
rect 425796 128460 425848 128512
rect 434628 128460 434680 128512
rect 419264 128392 419316 128444
rect 437480 128392 437532 128444
rect 141792 128324 141844 128376
rect 186320 128324 186372 128376
rect 412456 128324 412508 128376
rect 542360 128324 542412 128376
rect 131212 128256 131264 128308
rect 142804 128256 142856 128308
rect 131764 128188 131816 128240
rect 135996 128188 136048 128240
rect 411260 127032 411312 127084
rect 435456 127032 435508 127084
rect 140504 126964 140556 127016
rect 186320 126964 186372 127016
rect 413836 126964 413888 127016
rect 437480 126964 437532 127016
rect 131120 126896 131172 126948
rect 157984 126896 158036 126948
rect 131212 126828 131264 126880
rect 135904 126828 135956 126880
rect 131120 125672 131172 125724
rect 134524 125672 134576 125724
rect 144552 125604 144604 125656
rect 186320 125604 186372 125656
rect 413744 125604 413796 125656
rect 437480 125604 437532 125656
rect 131212 125536 131264 125588
rect 186964 125536 187016 125588
rect 131580 125468 131632 125520
rect 141424 125468 141476 125520
rect 411260 124244 411312 124296
rect 416228 124244 416280 124296
rect 141976 124176 142028 124228
rect 186320 124176 186372 124228
rect 413652 124176 413704 124228
rect 437480 124176 437532 124228
rect 131764 124108 131816 124160
rect 156604 124108 156656 124160
rect 131120 124040 131172 124092
rect 136088 124040 136140 124092
rect 411260 122884 411312 122936
rect 428556 122884 428608 122936
rect 144644 122816 144696 122868
rect 186320 122816 186372 122868
rect 413560 122816 413612 122868
rect 437480 122816 437532 122868
rect 131120 122748 131172 122800
rect 155224 122748 155276 122800
rect 131212 122680 131264 122732
rect 141516 122680 141568 122732
rect 131488 122612 131540 122664
rect 133236 122612 133288 122664
rect 423772 121524 423824 121576
rect 425796 121524 425848 121576
rect 141424 121456 141476 121508
rect 186320 121456 186372 121508
rect 131212 121388 131264 121440
rect 187056 121388 187108 121440
rect 131120 121320 131172 121372
rect 142896 121320 142948 121372
rect 410616 120708 410668 120760
rect 423772 120708 423824 120760
rect 411260 120096 411312 120148
rect 436836 120096 436888 120148
rect 131120 120028 131172 120080
rect 152464 120028 152516 120080
rect 132316 119960 132368 120012
rect 134616 119960 134668 120012
rect 142804 118668 142856 118720
rect 186320 118668 186372 118720
rect 411260 118668 411312 118720
rect 416320 118668 416372 118720
rect 131304 118600 131356 118652
rect 151084 118600 151136 118652
rect 131212 118532 131264 118584
rect 134708 118532 134760 118584
rect 131120 118464 131172 118516
rect 134800 118464 134852 118516
rect 134616 117376 134668 117428
rect 186412 117376 186464 117428
rect 131856 117308 131908 117360
rect 186320 117308 186372 117360
rect 131212 117240 131264 117292
rect 148324 117240 148376 117292
rect 131120 117172 131172 117224
rect 134892 117172 134944 117224
rect 142896 115948 142948 116000
rect 186320 115948 186372 116000
rect 132316 115880 132368 115932
rect 145564 115880 145616 115932
rect 131212 115472 131264 115524
rect 134984 115472 135036 115524
rect 134524 114520 134576 114572
rect 186320 114520 186372 114572
rect 411260 114520 411312 114572
rect 419172 114520 419224 114572
rect 131304 114452 131356 114504
rect 147036 114452 147088 114504
rect 411904 114452 411956 114504
rect 437480 114452 437532 114504
rect 131212 114384 131264 114436
rect 146944 114384 146996 114436
rect 131120 114316 131172 114368
rect 133328 114316 133380 114368
rect 131672 113160 131724 113212
rect 186320 113160 186372 113212
rect 411260 113160 411312 113212
rect 416412 113160 416464 113212
rect 131212 113092 131264 113144
rect 145656 113092 145708 113144
rect 412088 113092 412140 113144
rect 437480 113092 437532 113144
rect 131120 113024 131172 113076
rect 140136 113024 140188 113076
rect 135904 111868 135956 111920
rect 186412 111868 186464 111920
rect 134708 111800 134760 111852
rect 186320 111800 186372 111852
rect 131120 111732 131172 111784
rect 140044 111732 140096 111784
rect 131212 111664 131264 111716
rect 133420 111664 133472 111716
rect 131212 110372 131264 110424
rect 187148 110372 187200 110424
rect 421564 110372 421616 110424
rect 437480 110372 437532 110424
rect 131120 110304 131172 110356
rect 145748 110304 145800 110356
rect 131212 110236 131264 110288
rect 137284 110236 137336 110288
rect 135996 109012 136048 109064
rect 186320 109012 186372 109064
rect 411260 109012 411312 109064
rect 417976 109012 418028 109064
rect 131212 108944 131264 108996
rect 140228 108944 140280 108996
rect 416044 108944 416096 108996
rect 437480 108944 437532 108996
rect 131120 108876 131172 108928
rect 133604 108876 133656 108928
rect 131672 108468 131724 108520
rect 132316 108468 132368 108520
rect 131672 108332 131724 108384
rect 132040 108332 132092 108384
rect 131580 108264 131632 108316
rect 132132 108264 132184 108316
rect 133236 107652 133288 107704
rect 186320 107652 186372 107704
rect 411260 107652 411312 107704
rect 416504 107652 416556 107704
rect 131120 107584 131172 107636
rect 133512 107584 133564 107636
rect 411996 107584 412048 107636
rect 437480 107584 437532 107636
rect 131304 107516 131356 107568
rect 138664 107516 138716 107568
rect 131212 107448 131264 107500
rect 140320 107448 140372 107500
rect 140044 106292 140096 106344
rect 186320 106292 186372 106344
rect 131120 106224 131172 106276
rect 137376 106224 137428 106276
rect 131212 105952 131264 106004
rect 133696 105952 133748 106004
rect 136088 104932 136140 104984
rect 186412 104932 186464 104984
rect 134800 104864 134852 104916
rect 186320 104864 186372 104916
rect 131212 104796 131264 104848
rect 187240 104796 187292 104848
rect 421656 104796 421708 104848
rect 437480 104796 437532 104848
rect 131120 104728 131172 104780
rect 138756 104728 138808 104780
rect 411260 103504 411312 103556
rect 416044 103504 416096 103556
rect 131396 103436 131448 103488
rect 166264 103436 166316 103488
rect 131212 103368 131264 103420
rect 145840 103368 145892 103420
rect 131120 103300 131172 103352
rect 136180 103300 136232 103352
rect 435364 103028 435416 103080
rect 437664 103028 437716 103080
rect 134984 102144 135036 102196
rect 186320 102144 186372 102196
rect 131212 102076 131264 102128
rect 138848 102076 138900 102128
rect 416136 102076 416188 102128
rect 437480 102076 437532 102128
rect 134892 100716 134944 100768
rect 186320 100716 186372 100768
rect 411260 100716 411312 100768
rect 415124 100716 415176 100768
rect 131212 100648 131264 100700
rect 164884 100648 164936 100700
rect 432604 100648 432656 100700
rect 437480 100648 437532 100700
rect 540244 100648 540296 100700
rect 580172 100648 580224 100700
rect 131120 100580 131172 100632
rect 138940 100580 138992 100632
rect 140136 99424 140188 99476
rect 186412 99424 186464 99476
rect 136180 99356 136232 99408
rect 186320 99356 186372 99408
rect 131120 99288 131172 99340
rect 162124 99288 162176 99340
rect 131212 99220 131264 99272
rect 135076 99220 135128 99272
rect 133328 97996 133380 98048
rect 186320 97996 186372 98048
rect 131212 97928 131264 97980
rect 136272 97928 136324 97980
rect 431224 97928 431276 97980
rect 437480 97928 437532 97980
rect 140228 96636 140280 96688
rect 186320 96636 186372 96688
rect 131120 96568 131172 96620
rect 160744 96568 160796 96620
rect 429844 96568 429896 96620
rect 437480 96568 437532 96620
rect 131212 96500 131264 96552
rect 139032 96500 139084 96552
rect 131396 95888 131448 95940
rect 133788 95888 133840 95940
rect 411260 95820 411312 95872
rect 415216 95820 415268 95872
rect 144736 95208 144788 95260
rect 186320 95208 186372 95260
rect 131120 95140 131172 95192
rect 145932 95140 145984 95192
rect 428464 95140 428516 95192
rect 437480 95140 437532 95192
rect 131212 95072 131264 95124
rect 137468 95072 137520 95124
rect 411260 93916 411312 93968
rect 413376 93916 413428 93968
rect 133512 93848 133564 93900
rect 186320 93848 186372 93900
rect 131212 93780 131264 93832
rect 147128 93780 147180 93832
rect 425704 93780 425756 93832
rect 437480 93780 437532 93832
rect 131120 93712 131172 93764
rect 146024 93712 146076 93764
rect 138664 92556 138716 92608
rect 186412 92556 186464 92608
rect 131948 92488 132000 92540
rect 186320 92488 186372 92540
rect 131120 92420 131172 92472
rect 144184 92420 144236 92472
rect 411260 92420 411312 92472
rect 419356 92420 419408 92472
rect 424324 92420 424376 92472
rect 437480 92420 437532 92472
rect 131212 92352 131264 92404
rect 137560 92352 137612 92404
rect 133420 91060 133472 91112
rect 186320 91060 186372 91112
rect 132224 90992 132276 91044
rect 144276 90992 144328 91044
rect 421748 90992 421800 91044
rect 437480 90992 437532 91044
rect 131212 90924 131264 90976
rect 143080 90924 143132 90976
rect 411260 89768 411312 89820
rect 413376 89768 413428 89820
rect 138756 89700 138808 89752
rect 186320 89700 186372 89752
rect 131120 89632 131172 89684
rect 144368 89632 144420 89684
rect 418988 89632 419040 89684
rect 437480 89632 437532 89684
rect 131212 89564 131264 89616
rect 141608 89564 141660 89616
rect 132132 88340 132184 88392
rect 186320 88340 186372 88392
rect 131120 88272 131172 88324
rect 187332 88272 187384 88324
rect 411260 88272 411312 88324
rect 419264 88272 419316 88324
rect 420276 88272 420328 88324
rect 437480 88272 437532 88324
rect 131212 88204 131264 88256
rect 142988 88204 143040 88256
rect 131304 88136 131356 88188
rect 137652 88136 137704 88188
rect 133604 86980 133656 87032
rect 186320 86980 186372 87032
rect 131120 86912 131172 86964
rect 143172 86912 143224 86964
rect 131212 86844 131264 86896
rect 141700 86844 141752 86896
rect 411260 86436 411312 86488
rect 413836 86436 413888 86488
rect 131672 85552 131724 85604
rect 186320 85552 186372 85604
rect 131120 85484 131172 85536
rect 143264 85484 143316 85536
rect 417424 85484 417476 85536
rect 437480 85484 437532 85536
rect 131212 85416 131264 85468
rect 137744 85416 137796 85468
rect 142988 84192 143040 84244
rect 186320 84192 186372 84244
rect 131120 84124 131172 84176
rect 141884 84124 141936 84176
rect 411260 84124 411312 84176
rect 413744 84124 413796 84176
rect 420184 84124 420236 84176
rect 437480 84124 437532 84176
rect 131212 84056 131264 84108
rect 140412 84056 140464 84108
rect 131580 83988 131632 84040
rect 137836 83988 137888 84040
rect 131212 82764 131264 82816
rect 187424 82764 187476 82816
rect 417608 82764 417660 82816
rect 437480 82764 437532 82816
rect 131120 82696 131172 82748
rect 144460 82696 144512 82748
rect 132224 81404 132276 81456
rect 186320 81404 186372 81456
rect 411260 81404 411312 81456
rect 439504 81404 439556 81456
rect 131212 81336 131264 81388
rect 141792 81336 141844 81388
rect 420368 81336 420420 81388
rect 437480 81336 437532 81388
rect 131120 81268 131172 81320
rect 140504 81268 140556 81320
rect 133696 80044 133748 80096
rect 186320 80044 186372 80096
rect 131304 79976 131356 80028
rect 187516 79976 187568 80028
rect 417516 79976 417568 80028
rect 437480 79976 437532 80028
rect 131212 79908 131264 79960
rect 144552 79908 144604 79960
rect 131120 79840 131172 79892
rect 141976 79840 142028 79892
rect 131672 79296 131724 79348
rect 132040 79296 132092 79348
rect 135076 78684 135128 78736
rect 186320 78684 186372 78736
rect 131212 78616 131264 78668
rect 144644 78616 144696 78668
rect 419080 78616 419132 78668
rect 437480 78616 437532 78668
rect 131120 78548 131172 78600
rect 141424 78548 141476 78600
rect 411260 78208 411312 78260
rect 413652 78208 413704 78260
rect 141516 77256 141568 77308
rect 186320 77256 186372 77308
rect 417700 77188 417752 77240
rect 437480 77188 437532 77240
rect 131304 77120 131356 77172
rect 142804 77120 142856 77172
rect 131212 77052 131264 77104
rect 186964 77052 187016 77104
rect 411260 76712 411312 76764
rect 413468 76712 413520 76764
rect 131672 76576 131724 76628
rect 134616 76576 134668 76628
rect 131212 75828 131264 75880
rect 142896 75828 142948 75880
rect 134616 74604 134668 74656
rect 186412 74604 186464 74656
rect 133788 74536 133840 74588
rect 186320 74536 186372 74588
rect 131856 74468 131908 74520
rect 134524 74468 134576 74520
rect 414940 74468 414992 74520
rect 437480 74468 437532 74520
rect 411260 74196 411312 74248
rect 413560 74196 413612 74248
rect 131304 73108 131356 73160
rect 187056 73108 187108 73160
rect 411260 73108 411312 73160
rect 438492 73108 438544 73160
rect 131212 73040 131264 73092
rect 135904 73040 135956 73092
rect 417792 73040 417844 73092
rect 437480 73040 437532 73092
rect 131120 72972 131172 73024
rect 134708 72972 134760 73024
rect 151084 71748 151136 71800
rect 186320 71748 186372 71800
rect 131120 71680 131172 71732
rect 133236 71680 133288 71732
rect 415032 71680 415084 71732
rect 437480 71680 437532 71732
rect 131212 71612 131264 71664
rect 135996 71612 136048 71664
rect 134524 70388 134576 70440
rect 186320 70388 186372 70440
rect 131212 70320 131264 70372
rect 140044 70320 140096 70372
rect 421840 70320 421892 70372
rect 437480 70320 437532 70372
rect 131120 70252 131172 70304
rect 136088 70252 136140 70304
rect 131580 69640 131632 69692
rect 132040 69640 132092 69692
rect 137284 69096 137336 69148
rect 186320 69096 186372 69148
rect 131856 69028 131908 69080
rect 186412 69028 186464 69080
rect 411352 69028 411404 69080
rect 418988 69028 419040 69080
rect 131396 68960 131448 69012
rect 187148 68960 187200 69012
rect 411260 68960 411312 69012
rect 438400 68960 438452 69012
rect 131212 68892 131264 68944
rect 134800 68892 134852 68944
rect 417884 68892 417936 68944
rect 437480 68892 437532 68944
rect 131120 68824 131172 68876
rect 134984 68824 135036 68876
rect 148324 67600 148376 67652
rect 186320 67600 186372 67652
rect 131120 67532 131172 67584
rect 140136 67532 140188 67584
rect 429936 67532 429988 67584
rect 437480 67532 437532 67584
rect 131212 67328 131264 67380
rect 134892 67328 134944 67380
rect 133236 66240 133288 66292
rect 186320 66240 186372 66292
rect 411260 66240 411312 66292
rect 436744 66240 436796 66292
rect 131212 66172 131264 66224
rect 136180 66172 136232 66224
rect 421932 66172 421984 66224
rect 437480 66172 437532 66224
rect 131120 66104 131172 66156
rect 133328 66104 133380 66156
rect 132132 64880 132184 64932
rect 186320 64880 186372 64932
rect 131304 64812 131356 64864
rect 144736 64812 144788 64864
rect 431316 64812 431368 64864
rect 437480 64812 437532 64864
rect 131212 64744 131264 64796
rect 140228 64744 140280 64796
rect 131120 64676 131172 64728
rect 133512 64676 133564 64728
rect 411260 64472 411312 64524
rect 413284 64472 413336 64524
rect 146944 63520 146996 63572
rect 186320 63520 186372 63572
rect 131212 63452 131264 63504
rect 138664 63452 138716 63504
rect 411260 63452 411312 63504
rect 438308 63452 438360 63504
rect 132408 62092 132460 62144
rect 186320 62092 186372 62144
rect 131120 62024 131172 62076
rect 138756 62024 138808 62076
rect 422024 62024 422076 62076
rect 437480 62024 437532 62076
rect 131212 61956 131264 62008
rect 133420 61956 133472 62008
rect 144184 60732 144236 60784
rect 186320 60732 186372 60784
rect 131120 60664 131172 60716
rect 187240 60664 187292 60716
rect 432696 60664 432748 60716
rect 437480 60664 437532 60716
rect 544384 60664 544436 60716
rect 579804 60664 579856 60716
rect 131212 60596 131264 60648
rect 133604 60596 133656 60648
rect 411260 59372 411312 59424
rect 417424 59372 417476 59424
rect 131212 59304 131264 59356
rect 142988 59304 143040 59356
rect 420460 59304 420512 59356
rect 437480 59304 437532 59356
rect 131948 57944 132000 57996
rect 186320 57944 186372 57996
rect 411260 57944 411312 57996
rect 439596 57944 439648 57996
rect 131212 57876 131264 57928
rect 187332 57876 187384 57928
rect 412180 57876 412232 57928
rect 437480 57876 437532 57928
rect 131212 57332 131264 57384
rect 133696 57332 133748 57384
rect 133328 56584 133380 56636
rect 186320 56584 186372 56636
rect 131212 56516 131264 56568
rect 187424 56516 187476 56568
rect 420552 56516 420604 56568
rect 437480 56516 437532 56568
rect 131120 56448 131172 56500
rect 135076 56448 135128 56500
rect 132040 55224 132092 55276
rect 186320 55224 186372 55276
rect 131212 55156 131264 55208
rect 187516 55156 187568 55208
rect 132132 55088 132184 55140
rect 141516 55088 141568 55140
rect 435456 54680 435508 54732
rect 437756 54680 437808 54732
rect 411260 54000 411312 54052
rect 413468 54000 413520 54052
rect 133420 53796 133472 53848
rect 186320 53796 186372 53848
rect 131672 53728 131724 53780
rect 133788 53728 133840 53780
rect 416228 53728 416280 53780
rect 437480 53728 437532 53780
rect 131212 53660 131264 53712
rect 134616 53660 134668 53712
rect 131120 53592 131172 53644
rect 186964 53592 187016 53644
rect 411260 52504 411312 52556
rect 413284 52504 413336 52556
rect 132224 52368 132276 52420
rect 151084 52368 151136 52420
rect 428556 52368 428608 52420
rect 437480 52368 437532 52420
rect 131212 52300 131264 52352
rect 134524 52300 134576 52352
rect 132224 51076 132276 51128
rect 186320 51076 186372 51128
rect 132132 51008 132184 51060
rect 137284 51008 137336 51060
rect 133512 49716 133564 49768
rect 186320 49716 186372 49768
rect 131212 49648 131264 49700
rect 148324 49648 148376 49700
rect 131304 49580 131356 49632
rect 133236 49580 133288 49632
rect 131856 48288 131908 48340
rect 186320 48288 186372 48340
rect 411260 48288 411312 48340
rect 417516 48288 417568 48340
rect 131212 48220 131264 48272
rect 187148 48220 187200 48272
rect 416320 48220 416372 48272
rect 437480 48220 437532 48272
rect 132224 48152 132276 48204
rect 146944 48152 146996 48204
rect 132500 46928 132552 46980
rect 186320 46928 186372 46980
rect 131120 46860 131172 46912
rect 144184 46860 144236 46912
rect 412272 46860 412324 46912
rect 437480 46860 437532 46912
rect 131120 45500 131172 45552
rect 133328 45500 133380 45552
rect 419172 45500 419224 45552
rect 437480 45500 437532 45552
rect 131212 45432 131264 45484
rect 187056 45432 187108 45484
rect 131212 44072 131264 44124
rect 187240 44072 187292 44124
rect 416412 44072 416464 44124
rect 437480 44072 437532 44124
rect 131672 42848 131724 42900
rect 186412 42848 186464 42900
rect 131304 42780 131356 42832
rect 186320 42780 186372 42832
rect 131120 42712 131172 42764
rect 187332 42712 187384 42764
rect 411904 42712 411956 42764
rect 437480 42712 437532 42764
rect 131212 42644 131264 42696
rect 133420 42644 133472 42696
rect 411260 42644 411312 42696
rect 414848 42644 414900 42696
rect 131120 41352 131172 41404
rect 186964 41352 187016 41404
rect 417976 41352 418028 41404
rect 437480 41352 437532 41404
rect 131212 41284 131264 41336
rect 133512 41284 133564 41336
rect 411260 41012 411312 41064
rect 414756 41012 414808 41064
rect 411904 40672 411956 40724
rect 412180 40672 412232 40724
rect 411260 38836 411312 38888
rect 414664 38836 414716 38888
rect 131212 38564 131264 38616
rect 187148 38564 187200 38616
rect 416504 38564 416556 38616
rect 437480 38564 437532 38616
rect 131120 38496 131172 38548
rect 186596 38496 186648 38548
rect 132132 37340 132184 37392
rect 186412 37340 186464 37392
rect 132040 37272 132092 37324
rect 186320 37272 186372 37324
rect 131212 37204 131264 37256
rect 186504 37204 186556 37256
rect 411996 37204 412048 37256
rect 437480 37204 437532 37256
rect 411260 37136 411312 37188
rect 438216 37136 438268 37188
rect 132224 35912 132276 35964
rect 186320 35912 186372 35964
rect 131212 35844 131264 35896
rect 187240 35844 187292 35896
rect 416044 35844 416096 35896
rect 437480 35844 437532 35896
rect 131120 35776 131172 35828
rect 186964 35776 187016 35828
rect 411260 35776 411312 35828
rect 418896 35776 418948 35828
rect 415124 34416 415176 34468
rect 437480 34416 437532 34468
rect 131120 33124 131172 33176
rect 186320 33124 186372 33176
rect 131212 33056 131264 33108
rect 186412 33056 186464 33108
rect 411260 33056 411312 33108
rect 438124 33056 438176 33108
rect 412088 32988 412140 33040
rect 437480 32988 437532 33040
rect 131304 31832 131356 31884
rect 186320 31832 186372 31884
rect 131212 31764 131264 31816
rect 186412 31764 186464 31816
rect 412272 31696 412324 31748
rect 542636 31696 542688 31748
rect 412548 31628 412600 31680
rect 542544 31628 542596 31680
rect 412364 31560 412416 31612
rect 437480 31560 437532 31612
rect 131120 31016 131172 31068
rect 186320 31016 186372 31068
rect 186688 30268 186740 30320
rect 580172 30268 580224 30320
rect 411260 30200 411312 30252
rect 542728 30200 542780 30252
rect 411904 30132 411956 30184
rect 542360 30132 542412 30184
rect 412456 30064 412508 30116
rect 542452 30064 542504 30116
rect 188436 29452 188488 29504
rect 258908 29452 258960 29504
rect 188528 29384 188580 29436
rect 299572 29384 299624 29436
rect 130476 29316 130528 29368
rect 242992 29316 243044 29368
rect 417516 29316 417568 29368
rect 468760 29316 468812 29368
rect 201500 29248 201552 29300
rect 202512 29248 202564 29300
rect 410616 29248 410668 29300
rect 413468 29248 413520 29300
rect 485780 29248 485832 29300
rect 193220 29180 193272 29232
rect 194416 29180 194468 29232
rect 410524 29180 410576 29232
rect 452568 29180 452620 29232
rect 580356 29180 580408 29232
rect 130384 29112 130436 29164
rect 364708 29112 364760 29164
rect 444288 29112 444340 29164
rect 580264 29112 580316 29164
rect 226984 29044 227036 29096
rect 580448 29044 580500 29096
rect 210608 28976 210660 29028
rect 580540 28976 580592 29028
rect 130568 28908 130620 28960
rect 381084 28908 381136 28960
rect 413376 28908 413428 28960
rect 535460 28908 535512 28960
rect 130660 28840 130712 28892
rect 372988 28840 373040 28892
rect 418988 28840 419040 28892
rect 518992 28840 519044 28892
rect 188712 28772 188764 28824
rect 389180 28772 389232 28824
rect 439504 28772 439556 28824
rect 527180 28772 527232 28824
rect 188896 28704 188948 28756
rect 356612 28704 356664 28756
rect 417424 28704 417476 28756
rect 502340 28704 502392 28756
rect 188988 28636 189040 28688
rect 348516 28636 348568 28688
rect 436744 28636 436796 28688
rect 510620 28636 510672 28688
rect 182824 28568 182876 28620
rect 340420 28568 340472 28620
rect 413284 28568 413336 28620
rect 477500 28568 477552 28620
rect 188160 28500 188212 28552
rect 332140 28500 332192 28552
rect 439596 28500 439648 28552
rect 494152 28500 494204 28552
rect 188252 28432 188304 28484
rect 324412 28432 324464 28484
rect 188804 28364 188856 28416
rect 316132 28364 316184 28416
rect 189816 28296 189868 28348
rect 307760 28296 307812 28348
rect 188620 28228 188672 28280
rect 283380 28228 283432 28280
rect 189908 28160 189960 28212
rect 275100 28160 275152 28212
rect 189724 28092 189776 28144
rect 267004 28092 267056 28144
rect 188344 28024 188396 28076
rect 234620 28024 234672 28076
rect 79968 27548 80020 27600
rect 460480 27548 460532 27600
rect 418804 20612 418856 20664
rect 579988 20612 580040 20664
rect 218060 6808 218112 6860
rect 580172 6808 580224 6860
rect 2688 4088 2740 4140
rect 201500 4088 201552 4140
rect 1308 4020 1360 4072
rect 193220 4020 193272 4072
rect 1676 3680 1728 3732
rect 2688 3680 2740 3732
rect 572 3612 624 3664
rect 1308 3612 1360 3664
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 48226 334248 48282 334257
rect 48226 334183 48282 334192
rect 48134 333024 48190 333033
rect 48134 332959 48190 332968
rect 47950 331120 48006 331129
rect 47950 331055 48006 331064
rect 47858 328536 47914 328545
rect 47858 328471 47914 328480
rect 47766 327584 47822 327593
rect 47766 327519 47822 327528
rect 47674 305688 47730 305697
rect 47674 305623 47730 305632
rect 47688 254726 47716 305623
rect 47676 254720 47728 254726
rect 47676 254662 47728 254668
rect 47780 254658 47808 327519
rect 47768 254652 47820 254658
rect 47768 254594 47820 254600
rect 47872 254590 47900 328471
rect 47964 256018 47992 331055
rect 48042 325816 48098 325825
rect 48042 325751 48098 325760
rect 47952 256012 48004 256018
rect 47952 255954 48004 255960
rect 47860 254584 47912 254590
rect 47860 254526 47912 254532
rect 48056 250510 48084 325751
rect 48044 250504 48096 250510
rect 48044 250446 48096 250452
rect 48148 231810 48176 332959
rect 48136 231804 48188 231810
rect 48136 231746 48188 231752
rect 48240 131782 48268 334183
rect 208306 334112 208362 334121
rect 208306 334047 208362 334056
rect 49606 330122 49662 330131
rect 49606 330057 49662 330066
rect 49514 307274 49570 307283
rect 49514 307209 49570 307218
rect 49528 251870 49556 307209
rect 49620 256086 49648 330057
rect 208214 330032 208270 330041
rect 208214 329967 208270 329976
rect 208122 328536 208178 328545
rect 208122 328471 208178 328480
rect 208030 327448 208086 327457
rect 208030 327383 208086 327392
rect 207018 325816 207074 325825
rect 207018 325751 207074 325760
rect 207032 325718 207060 325751
rect 204260 325712 204312 325718
rect 204260 325654 204312 325660
rect 207020 325712 207072 325718
rect 207020 325654 207072 325660
rect 193220 306400 193272 306406
rect 193220 306342 193272 306348
rect 190460 305040 190512 305046
rect 190460 304982 190512 304988
rect 55862 299568 55918 299577
rect 55862 299503 55918 299512
rect 55876 298178 55904 299503
rect 103242 298208 103298 298217
rect 55220 298172 55272 298178
rect 55220 298114 55272 298120
rect 55864 298172 55916 298178
rect 103242 298143 103298 298152
rect 55864 298114 55916 298120
rect 49608 256080 49660 256086
rect 49608 256022 49660 256028
rect 49516 251864 49568 251870
rect 49516 251806 49568 251812
rect 48228 131776 48280 131782
rect 48228 131718 48280 131724
rect 1308 131232 1360 131238
rect 1308 131174 1360 131180
rect 55128 131232 55180 131238
rect 55232 131186 55260 298114
rect 65706 298072 65762 298081
rect 65706 298007 65762 298016
rect 67546 298072 67602 298081
rect 67546 298007 67602 298016
rect 67822 298072 67878 298081
rect 67822 298007 67878 298016
rect 69938 298072 69994 298081
rect 69938 298007 69994 298016
rect 70214 298072 70270 298081
rect 70214 298007 70270 298016
rect 71502 298072 71558 298081
rect 71502 298007 71558 298016
rect 73066 298072 73122 298081
rect 73066 298007 73122 298016
rect 74446 298072 74502 298081
rect 74446 298007 74502 298016
rect 75826 298072 75882 298081
rect 75826 298007 75882 298016
rect 76838 298072 76894 298081
rect 76838 298007 76894 298016
rect 77114 298072 77170 298081
rect 77114 298007 77170 298016
rect 78586 298072 78642 298081
rect 78586 298007 78642 298016
rect 79874 298072 79930 298081
rect 79874 298007 79930 298016
rect 81254 298072 81310 298081
rect 81254 298007 81310 298016
rect 81806 298072 81862 298081
rect 81806 298007 81862 298016
rect 82634 298072 82690 298081
rect 82634 298007 82690 298016
rect 84014 298072 84070 298081
rect 84014 298007 84070 298016
rect 85302 298072 85358 298081
rect 85302 298007 85358 298016
rect 86774 298072 86830 298081
rect 86774 298007 86830 298016
rect 88154 298072 88210 298081
rect 88154 298007 88210 298016
rect 89626 298072 89682 298081
rect 89626 298007 89682 298016
rect 90914 298072 90970 298081
rect 90914 298007 90970 298016
rect 92386 298072 92442 298081
rect 92386 298007 92442 298016
rect 93306 298072 93362 298081
rect 93306 298007 93362 298016
rect 93674 298072 93730 298081
rect 93674 298007 93730 298016
rect 95054 298072 95110 298081
rect 95054 298007 95110 298016
rect 96526 298072 96582 298081
rect 96526 298007 96582 298016
rect 96710 298072 96766 298081
rect 96710 298007 96766 298016
rect 97814 298072 97870 298081
rect 97814 298007 97870 298016
rect 99286 298072 99342 298081
rect 99286 298007 99342 298016
rect 100574 298072 100630 298081
rect 100574 298007 100630 298016
rect 101862 298072 101918 298081
rect 101862 298007 101918 298016
rect 65720 297294 65748 298007
rect 65708 297288 65760 297294
rect 65708 297230 65760 297236
rect 67560 252550 67588 298007
rect 67836 297226 67864 298007
rect 67824 297220 67876 297226
rect 67824 297162 67876 297168
rect 69952 297090 69980 298007
rect 70228 297158 70256 298007
rect 71516 297498 71544 298007
rect 71504 297492 71556 297498
rect 71504 297434 71556 297440
rect 70216 297152 70268 297158
rect 70216 297094 70268 297100
rect 69940 297084 69992 297090
rect 69940 297026 69992 297032
rect 67548 252544 67600 252550
rect 67548 252486 67600 252492
rect 73080 250578 73108 298007
rect 73068 250572 73120 250578
rect 73068 250514 73120 250520
rect 74460 229090 74488 298007
rect 75840 262886 75868 298007
rect 76852 297362 76880 298007
rect 76840 297356 76892 297362
rect 76840 297298 76892 297304
rect 75828 262880 75880 262886
rect 75828 262822 75880 262828
rect 77128 253230 77156 298007
rect 78494 297936 78550 297945
rect 78494 297871 78550 297880
rect 78508 257378 78536 297871
rect 78496 257372 78548 257378
rect 78496 257314 78548 257320
rect 77116 253224 77168 253230
rect 77116 253166 77168 253172
rect 78600 233238 78628 298007
rect 79782 297936 79838 297945
rect 79782 297871 79838 297880
rect 79796 297022 79824 297871
rect 79784 297016 79836 297022
rect 79784 296958 79836 296964
rect 79888 260234 79916 298007
rect 81268 262954 81296 298007
rect 81346 297936 81402 297945
rect 81346 297871 81402 297880
rect 81256 262948 81308 262954
rect 81256 262890 81308 262896
rect 81360 261526 81388 297871
rect 81820 297430 81848 298007
rect 81808 297424 81860 297430
rect 81808 297366 81860 297372
rect 81348 261520 81400 261526
rect 81348 261462 81400 261468
rect 79876 260228 79928 260234
rect 79876 260170 79928 260176
rect 78588 233232 78640 233238
rect 78588 233174 78640 233180
rect 82648 230450 82676 298007
rect 84028 252074 84056 298007
rect 84106 297936 84162 297945
rect 84106 297871 84162 297880
rect 84016 252068 84068 252074
rect 84016 252010 84068 252016
rect 82636 230444 82688 230450
rect 82636 230386 82688 230392
rect 74448 229084 74500 229090
rect 74448 229026 74500 229032
rect 55180 131180 55260 131186
rect 55128 131174 55260 131180
rect 1320 4078 1348 131174
rect 2688 131164 2740 131170
rect 2688 131106 2740 131112
rect 55140 131158 55260 131174
rect 2700 4146 2728 131106
rect 55140 129962 55168 131158
rect 84120 130422 84148 297871
rect 85316 130490 85344 298007
rect 85394 297936 85450 297945
rect 85394 297871 85450 297880
rect 86682 297936 86738 297945
rect 86682 297871 86738 297880
rect 85408 130626 85436 297871
rect 85486 297120 85542 297129
rect 85486 297055 85542 297064
rect 85500 130694 85528 297055
rect 86696 263022 86724 297871
rect 86684 263016 86736 263022
rect 86684 262958 86736 262964
rect 86788 237386 86816 298007
rect 86866 297800 86922 297809
rect 86866 297735 86922 297744
rect 86776 237380 86828 237386
rect 86776 237322 86828 237328
rect 85488 130688 85540 130694
rect 85488 130630 85540 130636
rect 85396 130620 85448 130626
rect 85396 130562 85448 130568
rect 86880 130558 86908 297735
rect 88168 251938 88196 298007
rect 88246 297936 88302 297945
rect 88246 297871 88302 297880
rect 89534 297936 89590 297945
rect 89534 297871 89590 297880
rect 88156 251932 88208 251938
rect 88156 251874 88208 251880
rect 88260 131986 88288 297871
rect 89548 238746 89576 297871
rect 89536 238740 89588 238746
rect 89536 238682 89588 238688
rect 89640 234598 89668 298007
rect 90928 257446 90956 298007
rect 91006 297936 91062 297945
rect 91006 297871 91062 297880
rect 92294 297936 92350 297945
rect 92294 297871 92350 297880
rect 90916 257440 90968 257446
rect 90916 257382 90968 257388
rect 91020 252006 91048 297871
rect 91008 252000 91060 252006
rect 91008 251942 91060 251948
rect 89628 234592 89680 234598
rect 89628 234534 89680 234540
rect 88248 131980 88300 131986
rect 88248 131922 88300 131928
rect 92308 131850 92336 297871
rect 92400 131918 92428 298007
rect 93320 296750 93348 298007
rect 93582 297936 93638 297945
rect 93582 297871 93638 297880
rect 93308 296744 93360 296750
rect 93308 296686 93360 296692
rect 93596 241466 93624 297871
rect 93688 256154 93716 298007
rect 93676 256148 93728 256154
rect 93676 256090 93728 256096
rect 93584 241460 93636 241466
rect 93584 241402 93636 241408
rect 95068 235958 95096 298007
rect 95146 297936 95202 297945
rect 95146 297871 95202 297880
rect 96434 297936 96490 297945
rect 96434 297871 96490 297880
rect 95160 297566 95188 297871
rect 95148 297560 95200 297566
rect 95148 297502 95200 297508
rect 96448 237318 96476 297871
rect 96436 237312 96488 237318
rect 96436 237254 96488 237260
rect 95056 235952 95108 235958
rect 95056 235894 95108 235900
rect 92388 131912 92440 131918
rect 92388 131854 92440 131860
rect 92296 131844 92348 131850
rect 92296 131786 92348 131792
rect 96540 130762 96568 298007
rect 96724 296818 96752 298007
rect 97722 297936 97778 297945
rect 97722 297871 97778 297880
rect 96712 296812 96764 296818
rect 96712 296754 96764 296760
rect 97736 132190 97764 297871
rect 97724 132184 97776 132190
rect 97724 132126 97776 132132
rect 97828 132054 97856 298007
rect 99194 297936 99250 297945
rect 99194 297871 99250 297880
rect 99208 263090 99236 297871
rect 99196 263084 99248 263090
rect 99196 263026 99248 263032
rect 99300 240106 99328 298007
rect 100588 260166 100616 298007
rect 100666 297936 100722 297945
rect 100666 297871 100722 297880
rect 100576 260160 100628 260166
rect 100576 260102 100628 260108
rect 99288 240100 99340 240106
rect 99288 240042 99340 240048
rect 100680 132258 100708 297871
rect 101876 245614 101904 298007
rect 102046 297936 102102 297945
rect 102046 297871 102102 297880
rect 101954 297800 102010 297809
rect 101954 297735 102010 297744
rect 101864 245608 101916 245614
rect 101864 245550 101916 245556
rect 101968 244254 101996 297735
rect 101956 244248 102008 244254
rect 101956 244190 102008 244196
rect 102060 242894 102088 297871
rect 103256 296886 103284 298143
rect 103334 298072 103390 298081
rect 103334 298007 103390 298016
rect 104806 298072 104862 298081
rect 104806 298007 104862 298016
rect 106186 298072 106242 298081
rect 106186 298007 106242 298016
rect 106738 298072 106794 298081
rect 106738 298007 106794 298016
rect 107474 298072 107530 298081
rect 107474 298007 107530 298016
rect 108946 298072 109002 298081
rect 108946 298007 109002 298016
rect 110326 298072 110382 298081
rect 110326 298007 110382 298016
rect 111706 298072 111762 298081
rect 111706 298007 111762 298016
rect 112994 298072 113050 298081
rect 112994 298007 113050 298016
rect 114466 298072 114522 298081
rect 114466 298007 114522 298016
rect 115846 298072 115902 298081
rect 115846 298007 115902 298016
rect 117226 298072 117282 298081
rect 117226 298007 117282 298016
rect 103244 296880 103296 296886
rect 103244 296822 103296 296828
rect 102048 242888 102100 242894
rect 102048 242830 102100 242836
rect 103348 132326 103376 298007
rect 104714 297936 104770 297945
rect 104714 297871 104770 297880
rect 104728 263158 104756 297871
rect 104716 263152 104768 263158
rect 104716 263094 104768 263100
rect 104820 261594 104848 298007
rect 106094 297936 106150 297945
rect 106094 297871 106150 297880
rect 104808 261588 104860 261594
rect 104808 261530 104860 261536
rect 106108 249762 106136 297871
rect 106096 249756 106148 249762
rect 106096 249698 106148 249704
rect 106200 242826 106228 298007
rect 106752 296954 106780 298007
rect 106740 296948 106792 296954
rect 106740 296890 106792 296896
rect 107488 250646 107516 298007
rect 108854 297936 108910 297945
rect 108854 297871 108910 297880
rect 107476 250640 107528 250646
rect 107476 250582 107528 250588
rect 108868 249694 108896 297871
rect 108856 249688 108908 249694
rect 108856 249630 108908 249636
rect 106188 242820 106240 242826
rect 106188 242762 106240 242768
rect 103336 132320 103388 132326
rect 103336 132262 103388 132268
rect 100668 132252 100720 132258
rect 100668 132194 100720 132200
rect 108960 132122 108988 298007
rect 110340 263226 110368 298007
rect 110328 263220 110380 263226
rect 110328 263162 110380 263168
rect 111720 252142 111748 298007
rect 111708 252136 111760 252142
rect 111708 252078 111760 252084
rect 113008 248402 113036 298007
rect 113086 297936 113142 297945
rect 113086 297871 113142 297880
rect 112996 248396 113048 248402
rect 112996 248338 113048 248344
rect 113100 247042 113128 297871
rect 114480 250782 114508 298007
rect 114468 250776 114520 250782
rect 114468 250718 114520 250724
rect 115860 250714 115888 298007
rect 117240 250850 117268 298007
rect 130384 297560 130436 297566
rect 130384 297502 130436 297508
rect 117228 250844 117280 250850
rect 117228 250786 117280 250792
rect 115848 250708 115900 250714
rect 115848 250650 115900 250656
rect 113088 247036 113140 247042
rect 113088 246978 113140 246984
rect 108948 132116 109000 132122
rect 108948 132058 109000 132064
rect 97816 132048 97868 132054
rect 97816 131990 97868 131996
rect 104900 131164 104952 131170
rect 104900 131106 104952 131112
rect 96528 130756 96580 130762
rect 96528 130698 96580 130704
rect 86868 130552 86920 130558
rect 86868 130494 86920 130500
rect 85304 130484 85356 130490
rect 85304 130426 85356 130432
rect 84108 130416 84160 130422
rect 84108 130358 84160 130364
rect 54978 129934 55168 129962
rect 104912 129948 104940 131106
rect 79980 27606 80008 30056
rect 130396 29170 130424 297502
rect 130476 297492 130528 297498
rect 130476 297434 130528 297440
rect 130488 29374 130516 297434
rect 188528 297424 188580 297430
rect 188528 297366 188580 297372
rect 188436 297356 188488 297362
rect 188436 297298 188488 297304
rect 188344 297288 188396 297294
rect 188344 297230 188396 297236
rect 147680 253224 147732 253230
rect 147680 253166 147732 253172
rect 147692 252210 147720 253166
rect 147680 252204 147732 252210
rect 147680 252146 147732 252152
rect 187240 249824 187292 249830
rect 187240 249766 187292 249772
rect 187252 244274 187280 249766
rect 187516 249756 187568 249762
rect 187516 249698 187568 249704
rect 187424 248464 187476 248470
rect 187528 248441 187556 249698
rect 187608 249688 187660 249694
rect 187608 249630 187660 249636
rect 187620 249529 187648 249630
rect 187606 249520 187662 249529
rect 187606 249455 187662 249464
rect 187424 248406 187476 248412
rect 187514 248432 187570 248441
rect 187332 247036 187384 247042
rect 187332 246978 187384 246984
rect 187344 246129 187372 246978
rect 187330 246120 187386 246129
rect 187330 246055 187386 246064
rect 187436 244934 187464 248406
rect 187514 248367 187570 248376
rect 187608 248396 187660 248402
rect 187608 248338 187660 248344
rect 187620 247353 187648 248338
rect 187606 247344 187662 247353
rect 187606 247279 187662 247288
rect 187608 245608 187660 245614
rect 187608 245550 187660 245556
rect 187620 245041 187648 245550
rect 187606 245032 187662 245041
rect 187606 244967 187662 244976
rect 187436 244906 187648 244934
rect 186320 244248 186372 244254
rect 187252 244246 187556 244274
rect 186320 244190 186372 244196
rect 186332 243953 186360 244190
rect 186318 243944 186374 243953
rect 186318 243879 186374 243888
rect 186412 242888 186464 242894
rect 186412 242830 186464 242836
rect 186320 242820 186372 242826
rect 186320 242762 186372 242768
rect 186332 242729 186360 242762
rect 186318 242720 186374 242729
rect 186318 242655 186374 242664
rect 186424 241641 186452 242830
rect 186410 241632 186466 241641
rect 186410 241567 186466 241576
rect 186320 241460 186372 241466
rect 186320 241402 186372 241408
rect 186332 240553 186360 241402
rect 186318 240544 186374 240553
rect 186318 240479 186374 240488
rect 186320 240100 186372 240106
rect 186320 240042 186372 240048
rect 186332 239465 186360 240042
rect 186318 239456 186374 239465
rect 186318 239391 186374 239400
rect 186320 238740 186372 238746
rect 186320 238682 186372 238688
rect 186332 238241 186360 238682
rect 186318 238232 186374 238241
rect 186318 238167 186374 238176
rect 186412 237380 186464 237386
rect 186412 237322 186464 237328
rect 186320 237312 186372 237318
rect 186320 237254 186372 237260
rect 186332 237153 186360 237254
rect 186318 237144 186374 237153
rect 186318 237079 186374 237088
rect 186424 236065 186452 237322
rect 186410 236056 186466 236065
rect 186410 235991 186466 236000
rect 186320 235952 186372 235958
rect 186320 235894 186372 235900
rect 186332 234841 186360 235894
rect 186318 234832 186374 234841
rect 186318 234767 186374 234776
rect 186320 234592 186372 234598
rect 186320 234534 186372 234540
rect 186332 233753 186360 234534
rect 186318 233744 186374 233753
rect 186318 233679 186374 233688
rect 186320 233232 186372 233238
rect 186320 233174 186372 233180
rect 186332 232665 186360 233174
rect 186318 232656 186374 232665
rect 186318 232591 186374 232600
rect 186320 231804 186372 231810
rect 186320 231746 186372 231752
rect 186332 231441 186360 231746
rect 186318 231432 186374 231441
rect 186318 231367 186374 231376
rect 186320 230444 186372 230450
rect 186320 230386 186372 230392
rect 186332 229265 186360 230386
rect 186318 229256 186374 229265
rect 186318 229191 186374 229200
rect 186320 229084 186372 229090
rect 186320 229026 186372 229032
rect 186332 228177 186360 229026
rect 186318 228168 186374 228177
rect 186318 228103 186374 228112
rect 186686 225720 186742 225729
rect 186686 225655 186742 225664
rect 186318 222320 186374 222329
rect 186318 222255 186374 222264
rect 186332 222222 186360 222255
rect 169024 222216 169076 222222
rect 169024 222158 169076 222164
rect 186320 222216 186372 222222
rect 186320 222158 186372 222164
rect 131856 220856 131908 220862
rect 131856 220798 131908 220804
rect 131672 132252 131724 132258
rect 131672 132194 131724 132200
rect 130568 132184 130620 132190
rect 130568 132126 130620 132132
rect 130476 29368 130528 29374
rect 130476 29310 130528 29316
rect 130384 29164 130436 29170
rect 130384 29106 130436 29112
rect 130580 28966 130608 132126
rect 130660 130756 130712 130762
rect 130660 130698 130712 130704
rect 130568 28960 130620 28966
rect 130568 28902 130620 28908
rect 130672 28898 130700 130698
rect 131120 129736 131172 129742
rect 131118 129704 131120 129713
rect 131172 129704 131174 129713
rect 131118 129639 131174 129648
rect 131212 129668 131264 129674
rect 131212 129610 131264 129616
rect 131224 128625 131252 129610
rect 131210 128616 131266 128625
rect 131210 128551 131266 128560
rect 131212 128308 131264 128314
rect 131212 128250 131264 128256
rect 131224 127401 131252 128250
rect 131210 127392 131266 127401
rect 131210 127327 131266 127336
rect 131120 126948 131172 126954
rect 131120 126890 131172 126896
rect 131132 126177 131160 126890
rect 131212 126880 131264 126886
rect 131210 126848 131212 126857
rect 131264 126848 131266 126857
rect 131210 126783 131266 126792
rect 131118 126168 131174 126177
rect 131118 126103 131174 126112
rect 131120 125724 131172 125730
rect 131120 125666 131172 125672
rect 131132 125633 131160 125666
rect 131118 125624 131174 125633
rect 131118 125559 131174 125568
rect 131212 125588 131264 125594
rect 131212 125530 131264 125536
rect 131224 124545 131252 125530
rect 131580 125520 131632 125526
rect 131580 125462 131632 125468
rect 131592 125089 131620 125462
rect 131578 125080 131634 125089
rect 131578 125015 131634 125024
rect 131210 124536 131266 124545
rect 131210 124471 131266 124480
rect 131120 124092 131172 124098
rect 131120 124034 131172 124040
rect 131132 123321 131160 124034
rect 131118 123312 131174 123321
rect 131118 123247 131174 123256
rect 131684 122834 131712 132194
rect 131868 129169 131896 220798
rect 159364 219496 159416 219502
rect 159364 219438 159416 219444
rect 135996 218068 136048 218074
rect 135996 218010 136048 218016
rect 135904 216708 135956 216714
rect 135904 216650 135956 216656
rect 134524 213988 134576 213994
rect 134524 213930 134576 213936
rect 133236 207052 133288 207058
rect 133236 206994 133288 207000
rect 131948 167068 132000 167074
rect 131948 167010 132000 167016
rect 131854 129160 131910 129169
rect 131854 129095 131910 129104
rect 131764 128240 131816 128246
rect 131764 128182 131816 128188
rect 131776 127945 131804 128182
rect 131762 127936 131818 127945
rect 131762 127871 131818 127880
rect 131764 124160 131816 124166
rect 131764 124102 131816 124108
rect 131776 123865 131804 124102
rect 131762 123856 131818 123865
rect 131762 123791 131818 123800
rect 131684 122806 131804 122834
rect 131120 122800 131172 122806
rect 131120 122742 131172 122748
rect 131210 122768 131266 122777
rect 131132 121553 131160 122742
rect 131210 122703 131212 122712
rect 131264 122703 131266 122712
rect 131212 122674 131264 122680
rect 131488 122664 131540 122670
rect 131488 122606 131540 122612
rect 131500 122097 131528 122606
rect 131486 122088 131542 122097
rect 131486 122023 131542 122032
rect 131118 121544 131174 121553
rect 131118 121479 131174 121488
rect 131212 121440 131264 121446
rect 131212 121382 131264 121388
rect 131120 121372 131172 121378
rect 131120 121314 131172 121320
rect 131132 120329 131160 121314
rect 131224 121009 131252 121382
rect 131210 121000 131266 121009
rect 131210 120935 131266 120944
rect 131118 120320 131174 120329
rect 131118 120255 131174 120264
rect 131120 120080 131172 120086
rect 131120 120022 131172 120028
rect 131132 119241 131160 120022
rect 131118 119232 131174 119241
rect 131118 119167 131174 119176
rect 131304 118652 131356 118658
rect 131304 118594 131356 118600
rect 131212 118584 131264 118590
rect 131210 118552 131212 118561
rect 131264 118552 131266 118561
rect 131120 118516 131172 118522
rect 131210 118487 131266 118496
rect 131120 118458 131172 118464
rect 131132 117473 131160 118458
rect 131316 118017 131344 118594
rect 131302 118008 131358 118017
rect 131302 117943 131358 117952
rect 131118 117464 131174 117473
rect 131118 117399 131174 117408
rect 131212 117292 131264 117298
rect 131212 117234 131264 117240
rect 131120 117224 131172 117230
rect 131120 117166 131172 117172
rect 131132 116249 131160 117166
rect 131224 116929 131252 117234
rect 131210 116920 131266 116929
rect 131210 116855 131266 116864
rect 131118 116240 131174 116249
rect 131118 116175 131174 116184
rect 131212 115524 131264 115530
rect 131212 115466 131264 115472
rect 131224 115161 131252 115466
rect 131210 115152 131266 115161
rect 131210 115087 131266 115096
rect 131304 114504 131356 114510
rect 131210 114472 131266 114481
rect 131304 114446 131356 114452
rect 131210 114407 131212 114416
rect 131264 114407 131266 114416
rect 131212 114378 131264 114384
rect 131120 114368 131172 114374
rect 131120 114310 131172 114316
rect 131132 113937 131160 114310
rect 131118 113928 131174 113937
rect 131118 113863 131174 113872
rect 131316 113393 131344 114446
rect 131302 113384 131358 113393
rect 131302 113319 131358 113328
rect 131672 113212 131724 113218
rect 131672 113154 131724 113160
rect 131212 113144 131264 113150
rect 131212 113086 131264 113092
rect 131120 113076 131172 113082
rect 131120 113018 131172 113024
rect 131132 112169 131160 113018
rect 131224 112849 131252 113086
rect 131210 112840 131266 112849
rect 131210 112775 131266 112784
rect 131118 112160 131174 112169
rect 131118 112095 131174 112104
rect 131120 111784 131172 111790
rect 131120 111726 131172 111732
rect 131132 111081 131160 111726
rect 131212 111716 131264 111722
rect 131212 111658 131264 111664
rect 131224 111625 131252 111658
rect 131210 111616 131266 111625
rect 131210 111551 131266 111560
rect 131118 111072 131174 111081
rect 131118 111007 131174 111016
rect 131212 110424 131264 110430
rect 131210 110392 131212 110401
rect 131264 110392 131266 110401
rect 131120 110356 131172 110362
rect 131210 110327 131266 110336
rect 131120 110298 131172 110304
rect 131132 109313 131160 110298
rect 131212 110288 131264 110294
rect 131212 110230 131264 110236
rect 131224 109857 131252 110230
rect 131210 109848 131266 109857
rect 131210 109783 131266 109792
rect 131118 109304 131174 109313
rect 131118 109239 131174 109248
rect 131212 108996 131264 109002
rect 131212 108938 131264 108944
rect 131120 108928 131172 108934
rect 131120 108870 131172 108876
rect 131132 108089 131160 108870
rect 131224 108633 131252 108938
rect 131210 108624 131266 108633
rect 131210 108559 131266 108568
rect 131684 108526 131712 113154
rect 131672 108520 131724 108526
rect 131672 108462 131724 108468
rect 131672 108384 131724 108390
rect 131672 108326 131724 108332
rect 131580 108316 131632 108322
rect 131580 108258 131632 108264
rect 131118 108080 131174 108089
rect 131118 108015 131174 108024
rect 131120 107636 131172 107642
rect 131120 107578 131172 107584
rect 131132 107001 131160 107578
rect 131304 107568 131356 107574
rect 131210 107536 131266 107545
rect 131304 107510 131356 107516
rect 131210 107471 131212 107480
rect 131264 107471 131266 107480
rect 131212 107442 131264 107448
rect 131118 106992 131174 107001
rect 131118 106927 131174 106936
rect 131316 106321 131344 107510
rect 131302 106312 131358 106321
rect 131120 106276 131172 106282
rect 131302 106247 131358 106256
rect 131120 106218 131172 106224
rect 131132 105233 131160 106218
rect 131212 106004 131264 106010
rect 131212 105946 131264 105952
rect 131224 105777 131252 105946
rect 131210 105768 131266 105777
rect 131210 105703 131266 105712
rect 131118 105224 131174 105233
rect 131118 105159 131174 105168
rect 131212 104848 131264 104854
rect 131212 104790 131264 104796
rect 131120 104780 131172 104786
rect 131120 104722 131172 104728
rect 131132 104009 131160 104722
rect 131224 104553 131252 104790
rect 131210 104544 131266 104553
rect 131210 104479 131266 104488
rect 131118 104000 131174 104009
rect 131118 103935 131174 103944
rect 131396 103488 131448 103494
rect 131210 103456 131266 103465
rect 131396 103430 131448 103436
rect 131210 103391 131212 103400
rect 131264 103391 131266 103400
rect 131212 103362 131264 103368
rect 131120 103352 131172 103358
rect 131120 103294 131172 103300
rect 131132 102241 131160 103294
rect 131408 102785 131436 103430
rect 131394 102776 131450 102785
rect 131394 102711 131450 102720
rect 131118 102232 131174 102241
rect 131118 102167 131174 102176
rect 131212 102128 131264 102134
rect 131212 102070 131264 102076
rect 131224 101153 131252 102070
rect 131210 101144 131266 101153
rect 131210 101079 131266 101088
rect 131212 100700 131264 100706
rect 131212 100642 131264 100648
rect 131120 100632 131172 100638
rect 131120 100574 131172 100580
rect 131132 99929 131160 100574
rect 131224 100473 131252 100642
rect 131210 100464 131266 100473
rect 131210 100399 131266 100408
rect 131118 99920 131174 99929
rect 131118 99855 131174 99864
rect 131120 99340 131172 99346
rect 131120 99282 131172 99288
rect 131132 98161 131160 99282
rect 131212 99272 131264 99278
rect 131212 99214 131264 99220
rect 131224 98705 131252 99214
rect 131210 98696 131266 98705
rect 131210 98631 131266 98640
rect 131118 98152 131174 98161
rect 131118 98087 131174 98096
rect 131212 97980 131264 97986
rect 131212 97922 131264 97928
rect 131224 97617 131252 97922
rect 131210 97608 131266 97617
rect 131210 97543 131266 97552
rect 131592 97073 131620 108258
rect 131684 99385 131712 108326
rect 131670 99376 131726 99385
rect 131670 99311 131726 99320
rect 131578 97064 131634 97073
rect 131578 96999 131634 97008
rect 131120 96620 131172 96626
rect 131120 96562 131172 96568
rect 131132 95849 131160 96562
rect 131212 96552 131264 96558
rect 131212 96494 131264 96500
rect 131224 96393 131252 96494
rect 131210 96384 131266 96393
rect 131210 96319 131266 96328
rect 131396 95940 131448 95946
rect 131396 95882 131448 95888
rect 131118 95840 131174 95849
rect 131118 95775 131174 95784
rect 131408 95305 131436 95882
rect 131394 95296 131450 95305
rect 131394 95231 131450 95240
rect 131120 95192 131172 95198
rect 131120 95134 131172 95140
rect 131132 94081 131160 95134
rect 131212 95124 131264 95130
rect 131212 95066 131264 95072
rect 131224 94625 131252 95066
rect 131210 94616 131266 94625
rect 131210 94551 131266 94560
rect 131118 94072 131174 94081
rect 131118 94007 131174 94016
rect 131212 93832 131264 93838
rect 131212 93774 131264 93780
rect 131120 93764 131172 93770
rect 131120 93706 131172 93712
rect 131132 92857 131160 93706
rect 131224 93537 131252 93774
rect 131210 93528 131266 93537
rect 131210 93463 131266 93472
rect 131118 92848 131174 92857
rect 131118 92783 131174 92792
rect 131120 92472 131172 92478
rect 131120 92414 131172 92420
rect 131132 91769 131160 92414
rect 131212 92404 131264 92410
rect 131212 92346 131264 92352
rect 131224 92313 131252 92346
rect 131210 92304 131266 92313
rect 131210 92239 131266 92248
rect 131118 91760 131174 91769
rect 131118 91695 131174 91704
rect 131212 90976 131264 90982
rect 131212 90918 131264 90924
rect 131224 90001 131252 90918
rect 131210 89992 131266 90001
rect 131210 89927 131266 89936
rect 131120 89684 131172 89690
rect 131120 89626 131172 89632
rect 131132 88777 131160 89626
rect 131212 89616 131264 89622
rect 131212 89558 131264 89564
rect 131224 89457 131252 89558
rect 131210 89448 131266 89457
rect 131210 89383 131266 89392
rect 131118 88768 131174 88777
rect 131118 88703 131174 88712
rect 131120 88324 131172 88330
rect 131120 88266 131172 88272
rect 131132 87689 131160 88266
rect 131212 88256 131264 88262
rect 131210 88224 131212 88233
rect 131264 88224 131266 88233
rect 131210 88159 131266 88168
rect 131304 88188 131356 88194
rect 131304 88130 131356 88136
rect 131118 87680 131174 87689
rect 131118 87615 131174 87624
rect 131316 87009 131344 88130
rect 131302 87000 131358 87009
rect 131120 86964 131172 86970
rect 131302 86935 131358 86944
rect 131120 86906 131172 86912
rect 131132 86465 131160 86906
rect 131212 86896 131264 86902
rect 131212 86838 131264 86844
rect 131118 86456 131174 86465
rect 131118 86391 131174 86400
rect 131224 85921 131252 86838
rect 131210 85912 131266 85921
rect 131210 85847 131266 85856
rect 131672 85604 131724 85610
rect 131672 85546 131724 85552
rect 131120 85536 131172 85542
rect 131120 85478 131172 85484
rect 131132 84697 131160 85478
rect 131212 85468 131264 85474
rect 131212 85410 131264 85416
rect 131224 85377 131252 85410
rect 131210 85368 131266 85377
rect 131210 85303 131266 85312
rect 131118 84688 131174 84697
rect 131118 84623 131174 84632
rect 131120 84176 131172 84182
rect 131120 84118 131172 84124
rect 131210 84144 131266 84153
rect 131132 82929 131160 84118
rect 131210 84079 131212 84088
rect 131264 84079 131266 84088
rect 131212 84050 131264 84056
rect 131580 84040 131632 84046
rect 131580 83982 131632 83988
rect 131592 83609 131620 83982
rect 131578 83600 131634 83609
rect 131578 83535 131634 83544
rect 131118 82920 131174 82929
rect 131118 82855 131174 82864
rect 131212 82816 131264 82822
rect 131212 82758 131264 82764
rect 131120 82748 131172 82754
rect 131120 82690 131172 82696
rect 131132 81841 131160 82690
rect 131224 82385 131252 82758
rect 131210 82376 131266 82385
rect 131210 82311 131266 82320
rect 131118 81832 131174 81841
rect 131118 81767 131174 81776
rect 131212 81388 131264 81394
rect 131212 81330 131264 81336
rect 131120 81320 131172 81326
rect 131120 81262 131172 81268
rect 131132 80617 131160 81262
rect 131224 81161 131252 81330
rect 131210 81152 131266 81161
rect 131210 81087 131266 81096
rect 131118 80608 131174 80617
rect 131118 80543 131174 80552
rect 131304 80028 131356 80034
rect 131304 79970 131356 79976
rect 131212 79960 131264 79966
rect 131210 79928 131212 79937
rect 131264 79928 131266 79937
rect 131120 79892 131172 79898
rect 131210 79863 131266 79872
rect 131120 79834 131172 79840
rect 131132 79529 131160 79834
rect 131118 79520 131174 79529
rect 131118 79455 131174 79464
rect 131316 78849 131344 79970
rect 131684 79354 131712 85546
rect 131672 79348 131724 79354
rect 131672 79290 131724 79296
rect 131302 78840 131358 78849
rect 131302 78775 131358 78784
rect 131212 78668 131264 78674
rect 131212 78610 131264 78616
rect 131120 78600 131172 78606
rect 131120 78542 131172 78548
rect 131132 77761 131160 78542
rect 131224 78305 131252 78610
rect 131210 78296 131266 78305
rect 131210 78231 131266 78240
rect 131118 77752 131174 77761
rect 131118 77687 131174 77696
rect 131304 77172 131356 77178
rect 131304 77114 131356 77120
rect 131212 77104 131264 77110
rect 131210 77072 131212 77081
rect 131264 77072 131266 77081
rect 131210 77007 131266 77016
rect 131316 76537 131344 77114
rect 131672 76628 131724 76634
rect 131672 76570 131724 76576
rect 131302 76528 131358 76537
rect 131302 76463 131358 76472
rect 131684 75993 131712 76570
rect 131670 75984 131726 75993
rect 131670 75919 131726 75928
rect 131212 75880 131264 75886
rect 131212 75822 131264 75828
rect 131224 74769 131252 75822
rect 131210 74760 131266 74769
rect 131210 74695 131266 74704
rect 131304 73160 131356 73166
rect 131304 73102 131356 73108
rect 131212 73092 131264 73098
rect 131212 73034 131264 73040
rect 131120 73024 131172 73030
rect 131224 73001 131252 73034
rect 131120 72966 131172 72972
rect 131210 72992 131266 73001
rect 131132 72457 131160 72966
rect 131210 72927 131266 72936
rect 131118 72448 131174 72457
rect 131118 72383 131174 72392
rect 131316 71913 131344 73102
rect 131302 71904 131358 71913
rect 131302 71839 131358 71848
rect 131120 71732 131172 71738
rect 131120 71674 131172 71680
rect 131132 70689 131160 71674
rect 131212 71664 131264 71670
rect 131212 71606 131264 71612
rect 131224 71233 131252 71606
rect 131210 71224 131266 71233
rect 131210 71159 131266 71168
rect 131118 70680 131174 70689
rect 131118 70615 131174 70624
rect 131212 70372 131264 70378
rect 131212 70314 131264 70320
rect 131120 70304 131172 70310
rect 131120 70246 131172 70252
rect 131132 69465 131160 70246
rect 131224 70145 131252 70314
rect 131210 70136 131266 70145
rect 131210 70071 131266 70080
rect 131580 69692 131632 69698
rect 131580 69634 131632 69640
rect 131118 69456 131174 69465
rect 131118 69391 131174 69400
rect 131396 69012 131448 69018
rect 131396 68954 131448 68960
rect 131212 68944 131264 68950
rect 131210 68912 131212 68921
rect 131264 68912 131266 68921
rect 131120 68876 131172 68882
rect 131210 68847 131266 68856
rect 131120 68818 131172 68824
rect 131132 67833 131160 68818
rect 131408 68377 131436 68954
rect 131394 68368 131450 68377
rect 131394 68303 131450 68312
rect 131118 67824 131174 67833
rect 131118 67759 131174 67768
rect 131120 67584 131172 67590
rect 131120 67526 131172 67532
rect 131132 66609 131160 67526
rect 131212 67380 131264 67386
rect 131212 67322 131264 67328
rect 131224 67153 131252 67322
rect 131210 67144 131266 67153
rect 131210 67079 131266 67088
rect 131118 66600 131174 66609
rect 131118 66535 131174 66544
rect 131212 66224 131264 66230
rect 131212 66166 131264 66172
rect 131120 66156 131172 66162
rect 131120 66098 131172 66104
rect 131132 65385 131160 66098
rect 131224 66065 131252 66166
rect 131210 66056 131266 66065
rect 131210 65991 131266 66000
rect 131118 65376 131174 65385
rect 131118 65311 131174 65320
rect 131304 64864 131356 64870
rect 131210 64832 131266 64841
rect 131304 64806 131356 64812
rect 131210 64767 131212 64776
rect 131264 64767 131266 64776
rect 131212 64738 131264 64744
rect 131120 64728 131172 64734
rect 131120 64670 131172 64676
rect 131132 63753 131160 64670
rect 131316 64297 131344 64806
rect 131302 64288 131358 64297
rect 131302 64223 131358 64232
rect 131118 63744 131174 63753
rect 131118 63679 131174 63688
rect 131212 63504 131264 63510
rect 131212 63446 131264 63452
rect 131224 63073 131252 63446
rect 131210 63064 131266 63073
rect 131210 62999 131266 63008
rect 131120 62076 131172 62082
rect 131120 62018 131172 62024
rect 131132 61305 131160 62018
rect 131212 62008 131264 62014
rect 131210 61976 131212 61985
rect 131264 61976 131266 61985
rect 131210 61911 131266 61920
rect 131118 61296 131174 61305
rect 131118 61231 131174 61240
rect 131120 60716 131172 60722
rect 131120 60658 131172 60664
rect 131132 59537 131160 60658
rect 131212 60648 131264 60654
rect 131212 60590 131264 60596
rect 131224 60217 131252 60590
rect 131210 60208 131266 60217
rect 131210 60143 131266 60152
rect 131118 59528 131174 59537
rect 131118 59463 131174 59472
rect 131212 59356 131264 59362
rect 131212 59298 131264 59304
rect 131224 58449 131252 59298
rect 131592 58993 131620 69634
rect 131578 58984 131634 58993
rect 131578 58919 131634 58928
rect 131210 58440 131266 58449
rect 131210 58375 131266 58384
rect 131212 57928 131264 57934
rect 131210 57896 131212 57905
rect 131264 57896 131266 57905
rect 131210 57831 131266 57840
rect 131212 57384 131264 57390
rect 131212 57326 131264 57332
rect 131224 56681 131252 57326
rect 131210 56672 131266 56681
rect 131210 56607 131266 56616
rect 131212 56568 131264 56574
rect 131212 56510 131264 56516
rect 131120 56500 131172 56506
rect 131120 56442 131172 56448
rect 131132 55457 131160 56442
rect 131224 56137 131252 56510
rect 131210 56128 131266 56137
rect 131210 56063 131266 56072
rect 131118 55448 131174 55457
rect 131118 55383 131174 55392
rect 131212 55208 131264 55214
rect 131212 55150 131264 55156
rect 131224 54369 131252 55150
rect 131210 54360 131266 54369
rect 131210 54295 131266 54304
rect 131672 53780 131724 53786
rect 131672 53722 131724 53728
rect 131212 53712 131264 53718
rect 131210 53680 131212 53689
rect 131264 53680 131266 53689
rect 131120 53644 131172 53650
rect 131210 53615 131266 53624
rect 131120 53586 131172 53592
rect 131132 52601 131160 53586
rect 131684 53145 131712 53722
rect 131670 53136 131726 53145
rect 131670 53071 131726 53080
rect 131118 52592 131174 52601
rect 131118 52527 131174 52536
rect 131212 52352 131264 52358
rect 131212 52294 131264 52300
rect 131224 51377 131252 52294
rect 131210 51368 131266 51377
rect 131210 51303 131266 51312
rect 131212 49700 131264 49706
rect 131212 49642 131264 49648
rect 131224 49609 131252 49642
rect 131304 49632 131356 49638
rect 131210 49600 131266 49609
rect 131304 49574 131356 49580
rect 131210 49535 131266 49544
rect 131316 49065 131344 49574
rect 131302 49056 131358 49065
rect 131302 48991 131358 49000
rect 131212 48272 131264 48278
rect 131212 48214 131264 48220
rect 131224 47297 131252 48214
rect 131210 47288 131266 47297
rect 131210 47223 131266 47232
rect 131120 46912 131172 46918
rect 131120 46854 131172 46860
rect 131132 46209 131160 46854
rect 131118 46200 131174 46209
rect 131118 46135 131174 46144
rect 131120 45552 131172 45558
rect 131120 45494 131172 45500
rect 131210 45520 131266 45529
rect 131132 44441 131160 45494
rect 131210 45455 131212 45464
rect 131264 45455 131266 45464
rect 131212 45426 131264 45432
rect 131118 44432 131174 44441
rect 131118 44367 131174 44376
rect 131212 44124 131264 44130
rect 131212 44066 131264 44072
rect 131224 43761 131252 44066
rect 131210 43752 131266 43761
rect 131210 43687 131266 43696
rect 131672 42900 131724 42906
rect 131672 42842 131724 42848
rect 131304 42832 131356 42838
rect 131304 42774 131356 42780
rect 131120 42764 131172 42770
rect 131120 42706 131172 42712
rect 131132 41993 131160 42706
rect 131212 42696 131264 42702
rect 131210 42664 131212 42673
rect 131264 42664 131266 42673
rect 131210 42599 131266 42608
rect 131118 41984 131174 41993
rect 131118 41919 131174 41928
rect 131120 41404 131172 41410
rect 131120 41346 131172 41352
rect 131132 40361 131160 41346
rect 131212 41336 131264 41342
rect 131212 41278 131264 41284
rect 131224 40905 131252 41278
rect 131210 40896 131266 40905
rect 131210 40831 131266 40840
rect 131118 40352 131174 40361
rect 131118 40287 131174 40296
rect 131212 38616 131264 38622
rect 131210 38584 131212 38593
rect 131264 38584 131266 38593
rect 131120 38548 131172 38554
rect 131210 38519 131266 38528
rect 131120 38490 131172 38496
rect 131132 37913 131160 38490
rect 131118 37904 131174 37913
rect 131118 37839 131174 37848
rect 131212 37256 131264 37262
rect 131212 37198 131264 37204
rect 131224 36145 131252 37198
rect 131316 36825 131344 42774
rect 131684 37369 131712 42842
rect 131670 37360 131726 37369
rect 131670 37295 131726 37304
rect 131302 36816 131358 36825
rect 131302 36751 131358 36760
rect 131210 36136 131266 36145
rect 131210 36071 131266 36080
rect 131212 35896 131264 35902
rect 131212 35838 131264 35844
rect 131120 35828 131172 35834
rect 131120 35770 131172 35776
rect 131132 35057 131160 35770
rect 131224 35601 131252 35838
rect 131210 35592 131266 35601
rect 131210 35527 131266 35536
rect 131118 35048 131174 35057
rect 131118 34983 131174 34992
rect 131120 33176 131172 33182
rect 131120 33118 131172 33124
rect 131132 32065 131160 33118
rect 131212 33108 131264 33114
rect 131212 33050 131264 33056
rect 131224 32745 131252 33050
rect 131210 32736 131266 32745
rect 131210 32671 131266 32680
rect 131118 32056 131174 32065
rect 131118 31991 131174 32000
rect 131304 31884 131356 31890
rect 131304 31826 131356 31832
rect 131212 31816 131264 31822
rect 131212 31758 131264 31764
rect 131224 31521 131252 31758
rect 131210 31512 131266 31521
rect 131210 31447 131266 31456
rect 131120 31068 131172 31074
rect 131120 31010 131172 31016
rect 131132 30433 131160 31010
rect 131316 30977 131344 31826
rect 131302 30968 131358 30977
rect 131302 30903 131358 30912
rect 131118 30424 131174 30433
rect 131118 30359 131174 30368
rect 130660 28892 130712 28898
rect 130660 28834 130712 28840
rect 131776 28801 131804 122806
rect 131856 117360 131908 117366
rect 131856 117302 131908 117308
rect 131868 75313 131896 117302
rect 131960 101697 131988 167010
rect 132040 162920 132092 162926
rect 132040 162862 132092 162868
rect 132052 108390 132080 162862
rect 132132 158772 132184 158778
rect 132132 158714 132184 158720
rect 132040 108384 132092 108390
rect 132040 108326 132092 108332
rect 132144 108322 132172 158714
rect 132224 147688 132276 147694
rect 132224 147630 132276 147636
rect 132132 108316 132184 108322
rect 132132 108258 132184 108264
rect 131946 101688 132002 101697
rect 131946 101623 132002 101632
rect 131948 92540 132000 92546
rect 131948 92482 132000 92488
rect 131854 75304 131910 75313
rect 131854 75239 131910 75248
rect 131856 74520 131908 74526
rect 131856 74462 131908 74468
rect 131868 74225 131896 74462
rect 131854 74216 131910 74225
rect 131854 74151 131910 74160
rect 131856 69080 131908 69086
rect 131856 69022 131908 69028
rect 131868 50289 131896 69022
rect 131960 62529 131988 92482
rect 132236 91225 132264 147630
rect 133144 132320 133196 132326
rect 133144 132262 133196 132268
rect 132316 120012 132368 120018
rect 132316 119954 132368 119960
rect 132328 119785 132356 119954
rect 132314 119776 132370 119785
rect 132314 119711 132370 119720
rect 132316 115932 132368 115938
rect 132316 115874 132368 115880
rect 132328 115705 132356 115874
rect 132314 115696 132370 115705
rect 132314 115631 132370 115640
rect 132316 108520 132368 108526
rect 132316 108462 132368 108468
rect 132222 91216 132278 91225
rect 132222 91151 132278 91160
rect 132224 91044 132276 91050
rect 132224 90986 132276 90992
rect 132236 90545 132264 90986
rect 132222 90536 132278 90545
rect 132222 90471 132278 90480
rect 132132 88392 132184 88398
rect 132132 88334 132184 88340
rect 132040 79348 132092 79354
rect 132040 79290 132092 79296
rect 132052 69698 132080 79290
rect 132040 69692 132092 69698
rect 132040 69634 132092 69640
rect 132144 66722 132172 88334
rect 132224 81456 132276 81462
rect 132224 81398 132276 81404
rect 132052 66694 132172 66722
rect 131946 62520 132002 62529
rect 131946 62455 132002 62464
rect 132052 60761 132080 66694
rect 132132 64932 132184 64938
rect 132132 64874 132184 64880
rect 132038 60752 132094 60761
rect 132038 60687 132094 60696
rect 131948 57996 132000 58002
rect 131948 57938 132000 57944
rect 131854 50280 131910 50289
rect 131854 50215 131910 50224
rect 131856 48340 131908 48346
rect 131856 48282 131908 48288
rect 131868 39681 131896 48282
rect 131960 44985 131988 57938
rect 132040 55276 132092 55282
rect 132040 55218 132092 55224
rect 131946 44976 132002 44985
rect 131946 44911 132002 44920
rect 132052 43217 132080 55218
rect 132144 55214 132172 64874
rect 132236 57225 132264 81398
rect 132328 77194 132356 108462
rect 132328 77166 132540 77194
rect 132512 76974 132540 77166
rect 132328 76946 132540 76974
rect 132328 73681 132356 76946
rect 132314 73672 132370 73681
rect 132314 73607 132370 73616
rect 132408 62144 132460 62150
rect 132408 62086 132460 62092
rect 132222 57216 132278 57225
rect 132222 57151 132278 57160
rect 132144 55186 132356 55214
rect 132132 55140 132184 55146
rect 132132 55082 132184 55088
rect 132144 54913 132172 55082
rect 132130 54904 132186 54913
rect 132130 54839 132186 54848
rect 132224 52420 132276 52426
rect 132224 52362 132276 52368
rect 132236 52057 132264 52362
rect 132222 52048 132278 52057
rect 132222 51983 132278 51992
rect 132224 51128 132276 51134
rect 132224 51070 132276 51076
rect 132132 51060 132184 51066
rect 132132 51002 132184 51008
rect 132144 50833 132172 51002
rect 132130 50824 132186 50833
rect 132130 50759 132186 50768
rect 132236 48314 132264 51070
rect 132328 48521 132356 55186
rect 132314 48512 132370 48521
rect 132314 48447 132370 48456
rect 132144 48286 132264 48314
rect 132420 48314 132448 62086
rect 132420 48286 132540 48314
rect 132038 43208 132094 43217
rect 132038 43143 132094 43152
rect 132144 41449 132172 48286
rect 132224 48204 132276 48210
rect 132224 48146 132276 48152
rect 132236 47841 132264 48146
rect 132222 47832 132278 47841
rect 132222 47767 132278 47776
rect 132512 47734 132540 48286
rect 132420 47706 132540 47734
rect 132420 46753 132448 47706
rect 132500 46980 132552 46986
rect 132500 46922 132552 46928
rect 132406 46744 132462 46753
rect 132406 46679 132462 46688
rect 132130 41440 132186 41449
rect 132130 41375 132186 41384
rect 131854 39672 131910 39681
rect 131854 39607 131910 39616
rect 132512 39137 132540 46922
rect 132498 39128 132554 39137
rect 132498 39063 132554 39072
rect 132132 37392 132184 37398
rect 132132 37334 132184 37340
rect 132040 37324 132092 37330
rect 132040 37266 132092 37272
rect 132052 33833 132080 37266
rect 132144 34513 132172 37334
rect 132224 35964 132276 35970
rect 132224 35906 132276 35912
rect 132130 34504 132186 34513
rect 132130 34439 132186 34448
rect 132038 33824 132094 33833
rect 132038 33759 132094 33768
rect 132236 33289 132264 35906
rect 132222 33280 132278 33289
rect 132222 33215 132278 33224
rect 133156 28937 133184 132262
rect 133248 122670 133276 206994
rect 133328 191888 133380 191894
rect 133328 191830 133380 191836
rect 133236 122664 133288 122670
rect 133236 122606 133288 122612
rect 133340 114374 133368 191830
rect 133420 186380 133472 186386
rect 133420 186322 133472 186328
rect 133328 114368 133380 114374
rect 133328 114310 133380 114316
rect 133432 111722 133460 186322
rect 133604 179444 133656 179450
rect 133604 179386 133656 179392
rect 133512 178084 133564 178090
rect 133512 178026 133564 178032
rect 133420 111716 133472 111722
rect 133420 111658 133472 111664
rect 133236 107704 133288 107710
rect 133236 107646 133288 107652
rect 133248 71738 133276 107646
rect 133524 107642 133552 178026
rect 133616 108934 133644 179386
rect 133696 175296 133748 175302
rect 133696 175238 133748 175244
rect 133604 108928 133656 108934
rect 133604 108870 133656 108876
rect 133512 107636 133564 107642
rect 133512 107578 133564 107584
rect 133708 106010 133736 175238
rect 133788 154624 133840 154630
rect 133788 154566 133840 154572
rect 133696 106004 133748 106010
rect 133696 105946 133748 105952
rect 133328 98048 133380 98054
rect 133328 97990 133380 97996
rect 133236 71732 133288 71738
rect 133236 71674 133288 71680
rect 133236 66292 133288 66298
rect 133236 66234 133288 66240
rect 133248 49638 133276 66234
rect 133340 66162 133368 97990
rect 133800 95946 133828 154566
rect 134536 125730 134564 213930
rect 134616 202904 134668 202910
rect 134616 202846 134668 202852
rect 134524 125724 134576 125730
rect 134524 125666 134576 125672
rect 134628 120018 134656 202846
rect 134708 200184 134760 200190
rect 134708 200126 134760 200132
rect 134616 120012 134668 120018
rect 134616 119954 134668 119960
rect 134720 118590 134748 200126
rect 134800 198756 134852 198762
rect 134800 198698 134852 198704
rect 134708 118584 134760 118590
rect 134708 118526 134760 118532
rect 134812 118522 134840 198698
rect 134892 196036 134944 196042
rect 134892 195978 134944 195984
rect 134800 118516 134852 118522
rect 134800 118458 134852 118464
rect 134616 117428 134668 117434
rect 134616 117370 134668 117376
rect 134524 114572 134576 114578
rect 134524 114514 134576 114520
rect 133788 95940 133840 95946
rect 133788 95882 133840 95888
rect 133512 93900 133564 93906
rect 133512 93842 133564 93848
rect 133420 91112 133472 91118
rect 133420 91054 133472 91060
rect 133328 66156 133380 66162
rect 133328 66098 133380 66104
rect 133432 62014 133460 91054
rect 133524 64734 133552 93842
rect 133604 87032 133656 87038
rect 133604 86974 133656 86980
rect 133512 64728 133564 64734
rect 133512 64670 133564 64676
rect 133420 62008 133472 62014
rect 133420 61950 133472 61956
rect 133616 60654 133644 86974
rect 133696 80096 133748 80102
rect 133696 80038 133748 80044
rect 133604 60648 133656 60654
rect 133604 60590 133656 60596
rect 133708 57390 133736 80038
rect 133788 74588 133840 74594
rect 133788 74530 133840 74536
rect 133696 57384 133748 57390
rect 133696 57326 133748 57332
rect 133328 56636 133380 56642
rect 133328 56578 133380 56584
rect 133236 49632 133288 49638
rect 133236 49574 133288 49580
rect 133340 45558 133368 56578
rect 133420 53848 133472 53854
rect 133420 53790 133472 53796
rect 133328 45552 133380 45558
rect 133328 45494 133380 45500
rect 133432 42702 133460 53790
rect 133800 53786 133828 74530
rect 134536 74526 134564 114514
rect 134628 76634 134656 117370
rect 134904 117230 134932 195978
rect 134984 193248 135036 193254
rect 134984 193190 135036 193196
rect 134892 117224 134944 117230
rect 134892 117166 134944 117172
rect 134996 115530 135024 193190
rect 135076 161492 135128 161498
rect 135076 161434 135128 161440
rect 134984 115524 135036 115530
rect 134984 115466 135036 115472
rect 134708 111852 134760 111858
rect 134708 111794 134760 111800
rect 134616 76628 134668 76634
rect 134616 76570 134668 76576
rect 134616 74656 134668 74662
rect 134616 74598 134668 74604
rect 134524 74520 134576 74526
rect 134524 74462 134576 74468
rect 134524 70440 134576 70446
rect 134524 70382 134576 70388
rect 133788 53780 133840 53786
rect 133788 53722 133840 53728
rect 134536 52358 134564 70382
rect 134628 53718 134656 74598
rect 134720 73030 134748 111794
rect 134800 104916 134852 104922
rect 134800 104858 134852 104864
rect 134708 73024 134760 73030
rect 134708 72966 134760 72972
rect 134812 68950 134840 104858
rect 134984 102196 135036 102202
rect 134984 102138 135036 102144
rect 134892 100768 134944 100774
rect 134892 100710 134944 100716
rect 134800 68944 134852 68950
rect 134800 68886 134852 68892
rect 134904 67386 134932 100710
rect 134996 68882 135024 102138
rect 135088 99278 135116 161434
rect 135916 126886 135944 216650
rect 136008 128246 136036 218010
rect 142804 216776 142856 216782
rect 142804 216718 142856 216724
rect 141424 212560 141476 212566
rect 141424 212502 141476 212508
rect 136088 209840 136140 209846
rect 136088 209782 136140 209788
rect 135996 128240 136048 128246
rect 135996 128182 136048 128188
rect 135904 126880 135956 126886
rect 135904 126822 135956 126828
rect 136100 124098 136128 209782
rect 140136 187740 140188 187746
rect 140136 187682 140188 187688
rect 140044 186448 140096 186454
rect 140044 186390 140096 186396
rect 137284 183592 137336 183598
rect 137284 183534 137336 183540
rect 136180 168428 136232 168434
rect 136180 168370 136232 168376
rect 136088 124092 136140 124098
rect 136088 124034 136140 124040
rect 135904 111920 135956 111926
rect 135904 111862 135956 111868
rect 135076 99272 135128 99278
rect 135076 99214 135128 99220
rect 135076 78736 135128 78742
rect 135076 78678 135128 78684
rect 134984 68876 135036 68882
rect 134984 68818 135036 68824
rect 134892 67380 134944 67386
rect 134892 67322 134944 67328
rect 135088 56506 135116 78678
rect 135916 73098 135944 111862
rect 135996 109064 136048 109070
rect 135996 109006 136048 109012
rect 135904 73092 135956 73098
rect 135904 73034 135956 73040
rect 136008 71670 136036 109006
rect 136088 104984 136140 104990
rect 136088 104926 136140 104932
rect 135996 71664 136048 71670
rect 135996 71606 136048 71612
rect 136100 70310 136128 104926
rect 136192 103358 136220 168370
rect 136272 160132 136324 160138
rect 136272 160074 136324 160080
rect 136180 103352 136232 103358
rect 136180 103294 136232 103300
rect 136180 99408 136232 99414
rect 136180 99350 136232 99356
rect 136088 70304 136140 70310
rect 136088 70246 136140 70252
rect 136192 66230 136220 99350
rect 136284 97986 136312 160074
rect 137296 110294 137324 183534
rect 138664 176724 138716 176730
rect 138664 176666 138716 176672
rect 137376 173936 137428 173942
rect 137376 173878 137428 173884
rect 137284 110288 137336 110294
rect 137284 110230 137336 110236
rect 137388 106282 137416 173878
rect 137468 154692 137520 154698
rect 137468 154634 137520 154640
rect 137376 106276 137428 106282
rect 137376 106218 137428 106224
rect 136272 97980 136324 97986
rect 136272 97922 136324 97928
rect 137480 95130 137508 154634
rect 137560 149116 137612 149122
rect 137560 149058 137612 149064
rect 137468 95124 137520 95130
rect 137468 95066 137520 95072
rect 137572 92410 137600 149058
rect 137652 139460 137704 139466
rect 137652 139402 137704 139408
rect 137560 92404 137612 92410
rect 137560 92346 137612 92352
rect 137664 88194 137692 139402
rect 137744 135312 137796 135318
rect 137744 135254 137796 135260
rect 137652 88188 137704 88194
rect 137652 88130 137704 88136
rect 137756 85474 137784 135254
rect 137836 132524 137888 132530
rect 137836 132466 137888 132472
rect 137744 85468 137796 85474
rect 137744 85410 137796 85416
rect 137848 84046 137876 132466
rect 138676 107574 138704 176666
rect 138756 172576 138808 172582
rect 138756 172518 138808 172524
rect 138664 107568 138716 107574
rect 138664 107510 138716 107516
rect 138768 104786 138796 172518
rect 138848 167136 138900 167142
rect 138848 167078 138900 167084
rect 138756 104780 138808 104786
rect 138756 104722 138808 104728
rect 138860 102134 138888 167078
rect 138940 164280 138992 164286
rect 138940 164222 138992 164228
rect 138848 102128 138900 102134
rect 138848 102070 138900 102076
rect 138952 100638 138980 164222
rect 139032 157412 139084 157418
rect 139032 157354 139084 157360
rect 138940 100632 138992 100638
rect 138940 100574 138992 100580
rect 139044 96558 139072 157354
rect 140056 111790 140084 186390
rect 140148 113082 140176 187682
rect 140228 180872 140280 180878
rect 140228 180814 140280 180820
rect 140136 113076 140188 113082
rect 140136 113018 140188 113024
rect 140044 111784 140096 111790
rect 140044 111726 140096 111732
rect 140240 109002 140268 180814
rect 140320 179512 140372 179518
rect 140320 179454 140372 179460
rect 140228 108996 140280 109002
rect 140228 108938 140280 108944
rect 140332 107506 140360 179454
rect 140412 133952 140464 133958
rect 140412 133894 140464 133900
rect 140320 107500 140372 107506
rect 140320 107442 140372 107448
rect 140044 106344 140096 106350
rect 140044 106286 140096 106292
rect 139032 96552 139084 96558
rect 139032 96494 139084 96500
rect 138664 92608 138716 92614
rect 138664 92550 138716 92556
rect 137836 84040 137888 84046
rect 137836 83982 137888 83988
rect 137284 69148 137336 69154
rect 137284 69090 137336 69096
rect 136180 66224 136232 66230
rect 136180 66166 136232 66172
rect 135076 56500 135128 56506
rect 135076 56442 135128 56448
rect 134616 53712 134668 53718
rect 134616 53654 134668 53660
rect 134524 52352 134576 52358
rect 134524 52294 134576 52300
rect 137296 51066 137324 69090
rect 138676 63510 138704 92550
rect 138756 89752 138808 89758
rect 138756 89694 138808 89700
rect 138664 63504 138716 63510
rect 138664 63446 138716 63452
rect 138768 62082 138796 89694
rect 140056 70378 140084 106286
rect 140136 99476 140188 99482
rect 140136 99418 140188 99424
rect 140044 70372 140096 70378
rect 140044 70314 140096 70320
rect 140148 67590 140176 99418
rect 140228 96688 140280 96694
rect 140228 96630 140280 96636
rect 140136 67584 140188 67590
rect 140136 67526 140188 67532
rect 140240 64802 140268 96630
rect 140424 84114 140452 133894
rect 140504 127016 140556 127022
rect 140504 126958 140556 126964
rect 140412 84108 140464 84114
rect 140412 84050 140464 84056
rect 140516 81326 140544 126958
rect 141436 125526 141464 212502
rect 141516 208412 141568 208418
rect 141516 208354 141568 208360
rect 141424 125520 141476 125526
rect 141424 125462 141476 125468
rect 141528 122738 141556 208354
rect 141608 143608 141660 143614
rect 141608 143550 141660 143556
rect 141516 122732 141568 122738
rect 141516 122674 141568 122680
rect 141424 121508 141476 121514
rect 141424 121450 141476 121456
rect 140504 81320 140556 81326
rect 140504 81262 140556 81268
rect 141436 78606 141464 121450
rect 141620 89622 141648 143550
rect 141700 136672 141752 136678
rect 141700 136614 141752 136620
rect 141608 89616 141660 89622
rect 141608 89558 141660 89564
rect 141712 86902 141740 136614
rect 141884 131164 141936 131170
rect 141884 131106 141936 131112
rect 141792 128376 141844 128382
rect 141792 128318 141844 128324
rect 141700 86896 141752 86902
rect 141700 86838 141752 86844
rect 141804 81394 141832 128318
rect 141896 84182 141924 131106
rect 142816 128314 142844 216718
rect 157984 215348 158036 215354
rect 157984 215290 158036 215296
rect 156604 211200 156656 211206
rect 156604 211142 156656 211148
rect 155224 205692 155276 205698
rect 155224 205634 155276 205640
rect 142896 204332 142948 204338
rect 142896 204274 142948 204280
rect 142804 128308 142856 128314
rect 142804 128250 142856 128256
rect 141976 124228 142028 124234
rect 141976 124170 142028 124176
rect 141884 84176 141936 84182
rect 141884 84118 141936 84124
rect 141792 81388 141844 81394
rect 141792 81330 141844 81336
rect 141988 79898 142016 124170
rect 142908 121378 142936 204274
rect 152464 201544 152516 201550
rect 152464 201486 152516 201492
rect 151084 198824 151136 198830
rect 151084 198766 151136 198772
rect 148324 197396 148376 197402
rect 148324 197338 148376 197344
rect 145564 194608 145616 194614
rect 145564 194550 145616 194556
rect 144184 149184 144236 149190
rect 144184 149126 144236 149132
rect 143080 144968 143132 144974
rect 143080 144910 143132 144916
rect 142988 142180 143040 142186
rect 142988 142122 143040 142128
rect 142896 121372 142948 121378
rect 142896 121314 142948 121320
rect 142804 118720 142856 118726
rect 142804 118662 142856 118668
rect 141976 79892 142028 79898
rect 141976 79834 142028 79840
rect 141424 78600 141476 78606
rect 141424 78542 141476 78548
rect 141516 77308 141568 77314
rect 141516 77250 141568 77256
rect 140228 64796 140280 64802
rect 140228 64738 140280 64744
rect 138756 62076 138808 62082
rect 138756 62018 138808 62024
rect 141528 55146 141556 77250
rect 142816 77178 142844 118662
rect 142896 116000 142948 116006
rect 142896 115942 142948 115948
rect 142804 77172 142856 77178
rect 142804 77114 142856 77120
rect 142908 75886 142936 115942
rect 143000 88262 143028 142122
rect 143092 90982 143120 144910
rect 143172 138032 143224 138038
rect 143172 137974 143224 137980
rect 143080 90976 143132 90982
rect 143080 90918 143132 90924
rect 142988 88256 143040 88262
rect 142988 88198 143040 88204
rect 143184 86970 143212 137974
rect 143264 135380 143316 135386
rect 143264 135322 143316 135328
rect 143172 86964 143224 86970
rect 143172 86906 143224 86912
rect 143276 85542 143304 135322
rect 144196 92478 144224 149126
rect 144276 146328 144328 146334
rect 144276 146270 144328 146276
rect 144184 92472 144236 92478
rect 144184 92414 144236 92420
rect 144288 91050 144316 146270
rect 144368 142248 144420 142254
rect 144368 142190 144420 142196
rect 144276 91044 144328 91050
rect 144276 90986 144328 90992
rect 144380 89690 144408 142190
rect 144460 129804 144512 129810
rect 144460 129746 144512 129752
rect 144368 89684 144420 89690
rect 144368 89626 144420 89632
rect 143264 85536 143316 85542
rect 143264 85478 143316 85484
rect 142988 84244 143040 84250
rect 142988 84186 143040 84192
rect 142896 75880 142948 75886
rect 142896 75822 142948 75828
rect 143000 59362 143028 84186
rect 144472 82754 144500 129746
rect 144552 125656 144604 125662
rect 144552 125598 144604 125604
rect 144460 82748 144512 82754
rect 144460 82690 144512 82696
rect 144564 79966 144592 125598
rect 144644 122868 144696 122874
rect 144644 122810 144696 122816
rect 144552 79960 144604 79966
rect 144552 79902 144604 79908
rect 144656 78674 144684 122810
rect 145576 115938 145604 194550
rect 146944 191956 146996 191962
rect 146944 191898 146996 191904
rect 145656 189100 145708 189106
rect 145656 189042 145708 189048
rect 145564 115932 145616 115938
rect 145564 115874 145616 115880
rect 145668 113150 145696 189042
rect 145748 182232 145800 182238
rect 145748 182174 145800 182180
rect 145656 113144 145708 113150
rect 145656 113086 145708 113092
rect 145760 110362 145788 182174
rect 145840 171148 145892 171154
rect 145840 171090 145892 171096
rect 145748 110356 145800 110362
rect 145748 110298 145800 110304
rect 145852 103426 145880 171090
rect 145932 153264 145984 153270
rect 145932 153206 145984 153212
rect 145840 103420 145892 103426
rect 145840 103362 145892 103368
rect 144736 95260 144788 95266
rect 144736 95202 144788 95208
rect 144644 78668 144696 78674
rect 144644 78610 144696 78616
rect 144748 64870 144776 95202
rect 145944 95198 145972 153206
rect 146024 150476 146076 150482
rect 146024 150418 146076 150424
rect 145932 95192 145984 95198
rect 145932 95134 145984 95140
rect 146036 93770 146064 150418
rect 146956 114442 146984 191898
rect 147036 190528 147088 190534
rect 147036 190470 147088 190476
rect 147048 114510 147076 190470
rect 147128 151836 147180 151842
rect 147128 151778 147180 151784
rect 147036 114504 147088 114510
rect 147036 114446 147088 114452
rect 146944 114436 146996 114442
rect 146944 114378 146996 114384
rect 147140 93838 147168 151778
rect 148336 117298 148364 197338
rect 151096 118658 151124 198766
rect 152476 120086 152504 201486
rect 155236 122806 155264 205634
rect 156616 124166 156644 211142
rect 157996 126954 158024 215290
rect 159376 129674 159404 219438
rect 166264 169788 166316 169794
rect 166264 169730 166316 169736
rect 164884 165640 164936 165646
rect 164884 165582 164936 165588
rect 162124 161560 162176 161566
rect 162124 161502 162176 161508
rect 160744 155984 160796 155990
rect 160744 155926 160796 155932
rect 159364 129668 159416 129674
rect 159364 129610 159416 129616
rect 157984 126948 158036 126954
rect 157984 126890 158036 126896
rect 156604 124160 156656 124166
rect 156604 124102 156656 124108
rect 155224 122800 155276 122806
rect 155224 122742 155276 122748
rect 152464 120080 152516 120086
rect 152464 120022 152516 120028
rect 151084 118652 151136 118658
rect 151084 118594 151136 118600
rect 148324 117292 148376 117298
rect 148324 117234 148376 117240
rect 160756 96626 160784 155926
rect 162136 99346 162164 161502
rect 164896 100706 164924 165582
rect 166276 103494 166304 169730
rect 169036 129742 169064 222158
rect 186318 221232 186374 221241
rect 186318 221167 186374 221176
rect 186332 220862 186360 221167
rect 186320 220856 186372 220862
rect 186320 220798 186372 220804
rect 186318 220008 186374 220017
rect 186318 219943 186374 219952
rect 186332 219502 186360 219943
rect 186320 219496 186372 219502
rect 186320 219438 186372 219444
rect 186318 218920 186374 218929
rect 186318 218855 186374 218864
rect 186332 218074 186360 218855
rect 186320 218068 186372 218074
rect 186320 218010 186372 218016
rect 186410 217832 186466 217841
rect 186410 217767 186466 217776
rect 186424 216782 186452 217767
rect 186412 216776 186464 216782
rect 186318 216744 186374 216753
rect 186412 216718 186464 216724
rect 186318 216679 186320 216688
rect 186372 216679 186374 216688
rect 186320 216650 186372 216656
rect 186318 215520 186374 215529
rect 186318 215455 186374 215464
rect 186332 215354 186360 215455
rect 186320 215348 186372 215354
rect 186320 215290 186372 215296
rect 186318 214432 186374 214441
rect 186318 214367 186374 214376
rect 186332 213994 186360 214367
rect 186320 213988 186372 213994
rect 186320 213930 186372 213936
rect 186318 213344 186374 213353
rect 186318 213279 186374 213288
rect 186332 212566 186360 213279
rect 186320 212560 186372 212566
rect 186320 212502 186372 212508
rect 186320 211200 186372 211206
rect 186318 211168 186320 211177
rect 186372 211168 186374 211177
rect 186318 211103 186374 211112
rect 186318 209944 186374 209953
rect 186318 209879 186374 209888
rect 186332 209846 186360 209879
rect 186320 209840 186372 209846
rect 186320 209782 186372 209788
rect 186318 208720 186374 208729
rect 186318 208655 186374 208664
rect 186332 208418 186360 208655
rect 186320 208412 186372 208418
rect 186320 208354 186372 208360
rect 186318 207632 186374 207641
rect 186318 207567 186374 207576
rect 186332 207058 186360 207567
rect 186320 207052 186372 207058
rect 186320 206994 186372 207000
rect 186318 206544 186374 206553
rect 186318 206479 186374 206488
rect 186332 205698 186360 206479
rect 186320 205692 186372 205698
rect 186320 205634 186372 205640
rect 186318 204368 186374 204377
rect 186318 204303 186320 204312
rect 186372 204303 186374 204312
rect 186320 204274 186372 204280
rect 186318 203144 186374 203153
rect 186318 203079 186374 203088
rect 186332 202910 186360 203079
rect 186320 202904 186372 202910
rect 186320 202846 186372 202852
rect 186318 202056 186374 202065
rect 186318 201991 186374 202000
rect 186332 201550 186360 201991
rect 186320 201544 186372 201550
rect 186320 201486 186372 201492
rect 186318 200832 186374 200841
rect 186318 200767 186374 200776
rect 186332 200190 186360 200767
rect 186320 200184 186372 200190
rect 186320 200126 186372 200132
rect 186410 199744 186466 199753
rect 186410 199679 186466 199688
rect 186424 198830 186452 199679
rect 186412 198824 186464 198830
rect 186318 198792 186374 198801
rect 186412 198766 186464 198772
rect 186318 198727 186320 198736
rect 186372 198727 186374 198736
rect 186320 198698 186372 198704
rect 186318 197568 186374 197577
rect 186318 197503 186374 197512
rect 186332 197402 186360 197503
rect 186320 197396 186372 197402
rect 186320 197338 186372 197344
rect 186318 196344 186374 196353
rect 186318 196279 186374 196288
rect 186332 196042 186360 196279
rect 186320 196036 186372 196042
rect 186320 195978 186372 195984
rect 186318 195256 186374 195265
rect 186318 195191 186374 195200
rect 186332 194614 186360 195191
rect 186320 194608 186372 194614
rect 186320 194550 186372 194556
rect 186318 194168 186374 194177
rect 186318 194103 186374 194112
rect 186332 193254 186360 194103
rect 186320 193248 186372 193254
rect 186320 193190 186372 193196
rect 186410 192944 186466 192953
rect 186410 192879 186466 192888
rect 186424 191962 186452 192879
rect 186412 191956 186464 191962
rect 186412 191898 186464 191904
rect 186320 191888 186372 191894
rect 186318 191856 186320 191865
rect 186372 191856 186374 191865
rect 186318 191791 186374 191800
rect 186318 190768 186374 190777
rect 186318 190703 186374 190712
rect 186332 190534 186360 190703
rect 186320 190528 186372 190534
rect 186320 190470 186372 190476
rect 186318 189544 186374 189553
rect 186318 189479 186374 189488
rect 186332 189106 186360 189479
rect 186320 189100 186372 189106
rect 186320 189042 186372 189048
rect 186318 188456 186374 188465
rect 186318 188391 186374 188400
rect 186332 187746 186360 188391
rect 186320 187740 186372 187746
rect 186320 187682 186372 187688
rect 186410 187368 186466 187377
rect 186410 187303 186466 187312
rect 186320 186448 186372 186454
rect 186318 186416 186320 186425
rect 186372 186416 186374 186425
rect 186424 186386 186452 187303
rect 186318 186351 186374 186360
rect 186412 186380 186464 186386
rect 186412 186322 186464 186328
rect 186318 183968 186374 183977
rect 186318 183903 186374 183912
rect 186332 183598 186360 183903
rect 186320 183592 186372 183598
rect 186320 183534 186372 183540
rect 186318 182880 186374 182889
rect 186318 182815 186374 182824
rect 186332 182238 186360 182815
rect 186320 182232 186372 182238
rect 186320 182174 186372 182180
rect 186318 181656 186374 181665
rect 186318 181591 186374 181600
rect 186332 180878 186360 181591
rect 186320 180872 186372 180878
rect 186320 180814 186372 180820
rect 186410 180568 186466 180577
rect 186410 180503 186466 180512
rect 186320 179512 186372 179518
rect 186318 179480 186320 179489
rect 186372 179480 186374 179489
rect 186424 179450 186452 180503
rect 186318 179415 186374 179424
rect 186412 179444 186464 179450
rect 186412 179386 186464 179392
rect 186318 178256 186374 178265
rect 186318 178191 186374 178200
rect 186332 178090 186360 178191
rect 186320 178084 186372 178090
rect 186320 178026 186372 178032
rect 186318 177168 186374 177177
rect 186318 177103 186374 177112
rect 186332 176730 186360 177103
rect 186320 176724 186372 176730
rect 186320 176666 186372 176672
rect 186318 176080 186374 176089
rect 186318 176015 186374 176024
rect 186332 175302 186360 176015
rect 186320 175296 186372 175302
rect 186320 175238 186372 175244
rect 186318 174992 186374 175001
rect 186318 174927 186374 174936
rect 186332 173942 186360 174927
rect 186320 173936 186372 173942
rect 186320 173878 186372 173884
rect 186318 172680 186374 172689
rect 186318 172615 186374 172624
rect 186332 172582 186360 172615
rect 186320 172576 186372 172582
rect 186320 172518 186372 172524
rect 186318 171592 186374 171601
rect 186318 171527 186374 171536
rect 186332 171154 186360 171527
rect 186320 171148 186372 171154
rect 186320 171090 186372 171096
rect 186318 170368 186374 170377
rect 186318 170303 186374 170312
rect 186332 169794 186360 170303
rect 186320 169788 186372 169794
rect 186320 169730 186372 169736
rect 186318 169280 186374 169289
rect 186318 169215 186374 169224
rect 186332 168434 186360 169215
rect 186320 168428 186372 168434
rect 186320 168370 186372 168376
rect 186410 168192 186466 168201
rect 186410 168127 186466 168136
rect 186320 167136 186372 167142
rect 186318 167104 186320 167113
rect 186372 167104 186374 167113
rect 186424 167074 186452 168127
rect 186318 167039 186374 167048
rect 186412 167068 186464 167074
rect 186412 167010 186464 167016
rect 186318 165880 186374 165889
rect 186318 165815 186374 165824
rect 186332 165646 186360 165815
rect 186320 165640 186372 165646
rect 186320 165582 186372 165588
rect 186318 164792 186374 164801
rect 186318 164727 186374 164736
rect 186332 164286 186360 164727
rect 186320 164280 186372 164286
rect 186320 164222 186372 164228
rect 186318 163704 186374 163713
rect 186318 163639 186374 163648
rect 186332 162926 186360 163639
rect 186320 162920 186372 162926
rect 186320 162862 186372 162868
rect 186410 162480 186466 162489
rect 186410 162415 186466 162424
rect 186320 161560 186372 161566
rect 186318 161528 186320 161537
rect 186372 161528 186374 161537
rect 186424 161498 186452 162415
rect 186318 161463 186374 161472
rect 186412 161492 186464 161498
rect 186412 161434 186464 161440
rect 186318 160304 186374 160313
rect 186318 160239 186374 160248
rect 186332 160138 186360 160239
rect 186320 160132 186372 160138
rect 186320 160074 186372 160080
rect 186318 159080 186374 159089
rect 186318 159015 186374 159024
rect 186332 158778 186360 159015
rect 186320 158772 186372 158778
rect 186320 158714 186372 158720
rect 186318 157992 186374 158001
rect 186318 157927 186374 157936
rect 186332 157418 186360 157927
rect 186320 157412 186372 157418
rect 186320 157354 186372 157360
rect 186318 156904 186374 156913
rect 186318 156839 186374 156848
rect 186332 155990 186360 156839
rect 186320 155984 186372 155990
rect 186320 155926 186372 155932
rect 186410 155816 186466 155825
rect 186410 155751 186466 155760
rect 186318 154728 186374 154737
rect 186318 154663 186320 154672
rect 186372 154663 186374 154672
rect 186320 154634 186372 154640
rect 186424 154630 186452 155751
rect 186412 154624 186464 154630
rect 186412 154566 186464 154572
rect 186318 153504 186374 153513
rect 186318 153439 186374 153448
rect 186332 153270 186360 153439
rect 186320 153264 186372 153270
rect 186320 153206 186372 153212
rect 186318 152416 186374 152425
rect 186318 152351 186374 152360
rect 186332 151842 186360 152351
rect 186320 151836 186372 151842
rect 186320 151778 186372 151784
rect 186318 151192 186374 151201
rect 186318 151127 186374 151136
rect 186332 150482 186360 151127
rect 186320 150476 186372 150482
rect 186320 150418 186372 150424
rect 186410 150104 186466 150113
rect 186410 150039 186466 150048
rect 186320 149184 186372 149190
rect 186318 149152 186320 149161
rect 186372 149152 186374 149161
rect 186424 149122 186452 150039
rect 186318 149087 186374 149096
rect 186412 149116 186464 149122
rect 186412 149058 186464 149064
rect 186318 147792 186374 147801
rect 186318 147727 186374 147736
rect 186332 147694 186360 147727
rect 186320 147688 186372 147694
rect 186320 147630 186372 147636
rect 186318 146704 186374 146713
rect 186318 146639 186374 146648
rect 186332 146334 186360 146639
rect 186320 146328 186372 146334
rect 186320 146270 186372 146276
rect 186318 145616 186374 145625
rect 186318 145551 186374 145560
rect 186332 144974 186360 145551
rect 186320 144968 186372 144974
rect 186320 144910 186372 144916
rect 186318 144528 186374 144537
rect 186318 144463 186374 144472
rect 186332 143614 186360 144463
rect 186320 143608 186372 143614
rect 186320 143550 186372 143556
rect 186410 143304 186466 143313
rect 186410 143239 186466 143248
rect 186424 142254 186452 143239
rect 186412 142248 186464 142254
rect 186318 142216 186374 142225
rect 186412 142190 186464 142196
rect 186318 142151 186320 142160
rect 186372 142151 186374 142160
rect 186320 142122 186372 142128
rect 186318 139904 186374 139913
rect 186318 139839 186374 139848
rect 186332 139466 186360 139839
rect 186320 139460 186372 139466
rect 186320 139402 186372 139408
rect 186318 138816 186374 138825
rect 186318 138751 186374 138760
rect 186332 138038 186360 138751
rect 186320 138032 186372 138038
rect 186320 137974 186372 137980
rect 186318 137728 186374 137737
rect 186318 137663 186374 137672
rect 186332 136678 186360 137663
rect 186320 136672 186372 136678
rect 186320 136614 186372 136620
rect 186410 136504 186466 136513
rect 186410 136439 186466 136448
rect 186318 135416 186374 135425
rect 186318 135351 186320 135360
rect 186372 135351 186374 135360
rect 186320 135322 186372 135328
rect 186424 135318 186452 136439
rect 186412 135312 186464 135318
rect 186412 135254 186464 135260
rect 186318 134328 186374 134337
rect 186318 134263 186374 134272
rect 186332 133958 186360 134263
rect 186320 133952 186372 133958
rect 186320 133894 186372 133900
rect 186318 133240 186374 133249
rect 186318 133175 186374 133184
rect 186332 132530 186360 133175
rect 186320 132524 186372 132530
rect 186320 132466 186372 132472
rect 186318 132016 186374 132025
rect 182824 131980 182876 131986
rect 186318 131951 186374 131960
rect 182824 131922 182876 131928
rect 169024 129736 169076 129742
rect 169024 129678 169076 129684
rect 166264 103488 166316 103494
rect 166264 103430 166316 103436
rect 164884 100700 164936 100706
rect 164884 100642 164936 100648
rect 162124 99340 162176 99346
rect 162124 99282 162176 99288
rect 160744 96620 160796 96626
rect 160744 96562 160796 96568
rect 147128 93832 147180 93838
rect 147128 93774 147180 93780
rect 146024 93764 146076 93770
rect 146024 93706 146076 93712
rect 151084 71800 151136 71806
rect 151084 71742 151136 71748
rect 148324 67652 148376 67658
rect 148324 67594 148376 67600
rect 144736 64864 144788 64870
rect 144736 64806 144788 64812
rect 146944 63572 146996 63578
rect 146944 63514 146996 63520
rect 144184 60784 144236 60790
rect 144184 60726 144236 60732
rect 142988 59356 143040 59362
rect 142988 59298 143040 59304
rect 141516 55140 141568 55146
rect 141516 55082 141568 55088
rect 137284 51060 137336 51066
rect 137284 51002 137336 51008
rect 133512 49768 133564 49774
rect 133512 49710 133564 49716
rect 133420 42696 133472 42702
rect 133420 42638 133472 42644
rect 133524 41342 133552 49710
rect 144196 46918 144224 60726
rect 146956 48210 146984 63514
rect 148336 49706 148364 67594
rect 151096 52426 151124 71742
rect 151084 52420 151136 52426
rect 151084 52362 151136 52368
rect 148324 49700 148376 49706
rect 148324 49642 148376 49648
rect 146944 48204 146996 48210
rect 146944 48146 146996 48152
rect 144184 46912 144236 46918
rect 144184 46854 144236 46860
rect 133512 41336 133564 41342
rect 133512 41278 133564 41284
rect 133142 28928 133198 28937
rect 133142 28863 133198 28872
rect 131762 28792 131818 28801
rect 131762 28727 131818 28736
rect 182836 28626 182864 131922
rect 186332 131170 186360 131951
rect 186320 131164 186372 131170
rect 186320 131106 186372 131112
rect 186318 129840 186374 129849
rect 186318 129775 186320 129784
rect 186372 129775 186374 129784
rect 186320 129746 186372 129752
rect 186318 128616 186374 128625
rect 186318 128551 186374 128560
rect 186332 128382 186360 128551
rect 186320 128376 186372 128382
rect 186320 128318 186372 128324
rect 186318 127528 186374 127537
rect 186318 127463 186374 127472
rect 186332 127022 186360 127463
rect 186320 127016 186372 127022
rect 186320 126958 186372 126964
rect 186318 126440 186374 126449
rect 186318 126375 186374 126384
rect 186332 125662 186360 126375
rect 186320 125656 186372 125662
rect 186320 125598 186372 125604
rect 186318 125216 186374 125225
rect 186318 125151 186374 125160
rect 186332 124234 186360 125151
rect 186320 124228 186372 124234
rect 186320 124170 186372 124176
rect 186318 123040 186374 123049
rect 186318 122975 186374 122984
rect 186332 122874 186360 122975
rect 186320 122868 186372 122874
rect 186320 122810 186372 122816
rect 186318 121952 186374 121961
rect 186318 121887 186374 121896
rect 186332 121514 186360 121887
rect 186320 121508 186372 121514
rect 186320 121450 186372 121456
rect 186318 119640 186374 119649
rect 186318 119575 186374 119584
rect 186332 118726 186360 119575
rect 186320 118720 186372 118726
rect 186320 118662 186372 118668
rect 186410 118552 186466 118561
rect 186410 118487 186466 118496
rect 186424 117434 186452 118487
rect 186412 117428 186464 117434
rect 186412 117370 186464 117376
rect 186320 117360 186372 117366
rect 186318 117328 186320 117337
rect 186372 117328 186374 117337
rect 186318 117263 186374 117272
rect 186318 116240 186374 116249
rect 186318 116175 186374 116184
rect 186332 116006 186360 116175
rect 186320 116000 186372 116006
rect 186320 115942 186372 115948
rect 186318 115152 186374 115161
rect 186318 115087 186374 115096
rect 186332 114578 186360 115087
rect 186320 114572 186372 114578
rect 186320 114514 186372 114520
rect 186318 114064 186374 114073
rect 186318 113999 186374 114008
rect 186332 113218 186360 113999
rect 186320 113212 186372 113218
rect 186320 113154 186372 113160
rect 186410 112840 186466 112849
rect 186410 112775 186466 112784
rect 186424 111926 186452 112775
rect 186412 111920 186464 111926
rect 186318 111888 186374 111897
rect 186412 111862 186464 111868
rect 186318 111823 186320 111832
rect 186372 111823 186374 111832
rect 186320 111794 186372 111800
rect 186318 109440 186374 109449
rect 186318 109375 186374 109384
rect 186332 109070 186360 109375
rect 186320 109064 186372 109070
rect 186320 109006 186372 109012
rect 186318 108352 186374 108361
rect 186318 108287 186374 108296
rect 186332 107710 186360 108287
rect 186320 107704 186372 107710
rect 186320 107646 186372 107652
rect 186318 107264 186374 107273
rect 186318 107199 186374 107208
rect 186332 106350 186360 107199
rect 186320 106344 186372 106350
rect 186320 106286 186372 106292
rect 186410 106040 186466 106049
rect 186410 105975 186466 105984
rect 186424 104990 186452 105975
rect 186412 104984 186464 104990
rect 186318 104952 186374 104961
rect 186412 104926 186464 104932
rect 186318 104887 186320 104896
rect 186372 104887 186374 104896
rect 186320 104858 186372 104864
rect 186318 102776 186374 102785
rect 186318 102711 186374 102720
rect 186332 102202 186360 102711
rect 186320 102196 186372 102202
rect 186320 102138 186372 102144
rect 186318 101552 186374 101561
rect 186318 101487 186374 101496
rect 186332 100774 186360 101487
rect 186320 100768 186372 100774
rect 186320 100710 186372 100716
rect 186410 100464 186466 100473
rect 186410 100399 186466 100408
rect 186318 99512 186374 99521
rect 186424 99482 186452 100399
rect 186318 99447 186374 99456
rect 186412 99476 186464 99482
rect 186332 99414 186360 99447
rect 186412 99418 186464 99424
rect 186320 99408 186372 99414
rect 186320 99350 186372 99356
rect 186318 98152 186374 98161
rect 186318 98087 186374 98096
rect 186332 98054 186360 98087
rect 186320 98048 186372 98054
rect 186320 97990 186372 97996
rect 186318 97064 186374 97073
rect 186318 96999 186374 97008
rect 186332 96694 186360 96999
rect 186320 96688 186372 96694
rect 186320 96630 186372 96636
rect 186318 95976 186374 95985
rect 186318 95911 186374 95920
rect 186332 95266 186360 95911
rect 186320 95260 186372 95266
rect 186320 95202 186372 95208
rect 186318 94752 186374 94761
rect 186318 94687 186374 94696
rect 186332 93906 186360 94687
rect 186320 93900 186372 93906
rect 186320 93842 186372 93848
rect 186410 93664 186466 93673
rect 186410 93599 186466 93608
rect 186424 92614 186452 93599
rect 186412 92608 186464 92614
rect 186318 92576 186374 92585
rect 186412 92550 186464 92556
rect 186318 92511 186320 92520
rect 186372 92511 186374 92520
rect 186320 92482 186372 92488
rect 186318 91488 186374 91497
rect 186318 91423 186374 91432
rect 186332 91118 186360 91423
rect 186320 91112 186372 91118
rect 186320 91054 186372 91060
rect 186318 90264 186374 90273
rect 186318 90199 186374 90208
rect 186332 89758 186360 90199
rect 186320 89752 186372 89758
rect 186320 89694 186372 89700
rect 186318 89176 186374 89185
rect 186318 89111 186374 89120
rect 186332 88398 186360 89111
rect 186320 88392 186372 88398
rect 186320 88334 186372 88340
rect 186318 88088 186374 88097
rect 186318 88023 186374 88032
rect 186332 87038 186360 88023
rect 186320 87032 186372 87038
rect 186320 86974 186372 86980
rect 186318 85776 186374 85785
rect 186318 85711 186374 85720
rect 186332 85610 186360 85711
rect 186320 85604 186372 85610
rect 186320 85546 186372 85552
rect 186318 84688 186374 84697
rect 186318 84623 186374 84632
rect 186332 84250 186360 84623
rect 186320 84244 186372 84250
rect 186320 84186 186372 84192
rect 186318 82376 186374 82385
rect 186318 82311 186374 82320
rect 186332 81462 186360 82311
rect 186320 81456 186372 81462
rect 186320 81398 186372 81404
rect 186318 81288 186374 81297
rect 186318 81223 186374 81232
rect 186332 80102 186360 81223
rect 186320 80096 186372 80102
rect 186320 80038 186372 80044
rect 186318 78976 186374 78985
rect 186318 78911 186374 78920
rect 186332 78742 186360 78911
rect 186320 78736 186372 78742
rect 186320 78678 186372 78684
rect 186318 77888 186374 77897
rect 186318 77823 186374 77832
rect 186332 77314 186360 77823
rect 186320 77308 186372 77314
rect 186320 77250 186372 77256
rect 186410 75576 186466 75585
rect 186410 75511 186466 75520
rect 186424 74662 186452 75511
rect 186412 74656 186464 74662
rect 186318 74624 186374 74633
rect 186412 74598 186464 74604
rect 186318 74559 186320 74568
rect 186372 74559 186374 74568
rect 186320 74530 186372 74536
rect 186318 72312 186374 72321
rect 186318 72247 186374 72256
rect 186332 71806 186360 72247
rect 186320 71800 186372 71806
rect 186320 71742 186372 71748
rect 186318 71088 186374 71097
rect 186318 71023 186374 71032
rect 186332 70446 186360 71023
rect 186320 70440 186372 70446
rect 186320 70382 186372 70388
rect 186318 70000 186374 70009
rect 186318 69935 186374 69944
rect 186332 69154 186360 69935
rect 186320 69148 186372 69154
rect 186320 69090 186372 69096
rect 186412 69080 186464 69086
rect 186410 69048 186412 69057
rect 186464 69048 186466 69057
rect 186410 68983 186466 68992
rect 186318 67688 186374 67697
rect 186318 67623 186320 67632
rect 186372 67623 186374 67632
rect 186320 67594 186372 67600
rect 186318 66600 186374 66609
rect 186318 66535 186374 66544
rect 186332 66298 186360 66535
rect 186320 66292 186372 66298
rect 186320 66234 186372 66240
rect 186318 65512 186374 65521
rect 186318 65447 186374 65456
rect 186332 64938 186360 65447
rect 186320 64932 186372 64938
rect 186320 64874 186372 64880
rect 186318 64288 186374 64297
rect 186318 64223 186374 64232
rect 186332 63578 186360 64223
rect 186320 63572 186372 63578
rect 186320 63514 186372 63520
rect 186318 62248 186374 62257
rect 186318 62183 186374 62192
rect 186332 62150 186360 62183
rect 186320 62144 186372 62150
rect 186320 62086 186372 62092
rect 186318 61024 186374 61033
rect 186318 60959 186374 60968
rect 186332 60790 186360 60959
rect 186320 60784 186372 60790
rect 186320 60726 186372 60732
rect 186318 58712 186374 58721
rect 186318 58647 186374 58656
rect 186332 58002 186360 58647
rect 186320 57996 186372 58002
rect 186320 57938 186372 57944
rect 186318 57624 186374 57633
rect 186318 57559 186374 57568
rect 186332 56642 186360 57559
rect 186320 56636 186372 56642
rect 186320 56578 186372 56584
rect 186318 55312 186374 55321
rect 186318 55247 186320 55256
rect 186372 55247 186374 55256
rect 186320 55218 186372 55224
rect 186318 54224 186374 54233
rect 186318 54159 186374 54168
rect 186332 53854 186360 54159
rect 186320 53848 186372 53854
rect 186320 53790 186372 53796
rect 186318 51912 186374 51921
rect 186318 51847 186374 51856
rect 186332 51134 186360 51847
rect 186320 51128 186372 51134
rect 186320 51070 186372 51076
rect 186318 50824 186374 50833
rect 186318 50759 186374 50768
rect 186332 49774 186360 50759
rect 186320 49768 186372 49774
rect 186320 49710 186372 49716
rect 186318 48512 186374 48521
rect 186318 48447 186374 48456
rect 186332 48346 186360 48447
rect 186320 48340 186372 48346
rect 186320 48282 186372 48288
rect 186318 47424 186374 47433
rect 186318 47359 186374 47368
rect 186332 46986 186360 47359
rect 186320 46980 186372 46986
rect 186320 46922 186372 46928
rect 186594 45112 186650 45121
rect 186594 45047 186650 45056
rect 186410 44024 186466 44033
rect 186410 43959 186466 43968
rect 186318 42936 186374 42945
rect 186424 42906 186452 43959
rect 186318 42871 186374 42880
rect 186412 42900 186464 42906
rect 186332 42838 186360 42871
rect 186412 42842 186464 42848
rect 186320 42832 186372 42838
rect 186320 42774 186372 42780
rect 186502 41712 186558 41721
rect 186502 41647 186558 41656
rect 186410 38448 186466 38457
rect 186410 38383 186466 38392
rect 186424 37398 186452 38383
rect 186412 37392 186464 37398
rect 186318 37360 186374 37369
rect 186412 37334 186464 37340
rect 186318 37295 186320 37304
rect 186372 37295 186374 37304
rect 186320 37266 186372 37272
rect 186516 37262 186544 41647
rect 186608 38554 186636 45047
rect 186596 38548 186648 38554
rect 186596 38490 186648 38496
rect 186504 37256 186556 37262
rect 186504 37198 186556 37204
rect 186318 36136 186374 36145
rect 186318 36071 186374 36080
rect 186332 35970 186360 36071
rect 186320 35964 186372 35970
rect 186320 35906 186372 35912
rect 186410 35048 186466 35057
rect 186410 34983 186466 34992
rect 186318 33824 186374 33833
rect 186318 33759 186374 33768
rect 186332 33182 186360 33759
rect 186320 33176 186372 33182
rect 186320 33118 186372 33124
rect 186424 33114 186452 34983
rect 186412 33108 186464 33114
rect 186412 33050 186464 33056
rect 186410 32736 186466 32745
rect 186410 32671 186466 32680
rect 186320 31884 186372 31890
rect 186320 31826 186372 31832
rect 186332 31793 186360 31826
rect 186424 31822 186452 32671
rect 186412 31816 186464 31822
rect 186318 31784 186374 31793
rect 186412 31758 186464 31764
rect 186318 31719 186374 31728
rect 186320 31068 186372 31074
rect 186320 31010 186372 31016
rect 186332 30569 186360 31010
rect 186318 30560 186374 30569
rect 186318 30495 186374 30504
rect 186700 30326 186728 225655
rect 187528 224777 187556 244246
rect 187514 224768 187570 224777
rect 187514 224703 187570 224712
rect 187620 223553 187648 244906
rect 187606 223544 187662 223553
rect 187606 223479 187662 223488
rect 186962 212120 187018 212129
rect 186962 212055 187018 212064
rect 186976 125594 187004 212055
rect 187054 205456 187110 205465
rect 187054 205391 187110 205400
rect 186964 125588 187016 125594
rect 186964 125530 187016 125536
rect 187068 121446 187096 205391
rect 187146 185056 187202 185065
rect 187146 184991 187202 185000
rect 187056 121440 187108 121446
rect 187056 121382 187108 121388
rect 186962 120728 187018 120737
rect 186962 120663 187018 120672
rect 186976 77110 187004 120663
rect 187054 110664 187110 110673
rect 187054 110599 187110 110608
rect 186964 77104 187016 77110
rect 186964 77046 187016 77052
rect 186962 73400 187018 73409
rect 186962 73335 187018 73344
rect 186976 53650 187004 73335
rect 187068 73166 187096 110599
rect 187160 110430 187188 184991
rect 187238 173768 187294 173777
rect 187238 173703 187294 173712
rect 187148 110424 187200 110430
rect 187148 110366 187200 110372
rect 187252 104854 187280 173703
rect 187330 141128 187386 141137
rect 187330 141063 187386 141072
rect 187240 104848 187292 104854
rect 187240 104790 187292 104796
rect 187146 103864 187202 103873
rect 187146 103799 187202 103808
rect 187056 73160 187108 73166
rect 187056 73102 187108 73108
rect 187160 69018 187188 103799
rect 187344 88330 187372 141063
rect 187422 130928 187478 130937
rect 187422 130863 187478 130872
rect 187332 88324 187384 88330
rect 187332 88266 187384 88272
rect 187238 87000 187294 87009
rect 187238 86935 187294 86944
rect 187148 69012 187200 69018
rect 187148 68954 187200 68960
rect 187146 63200 187202 63209
rect 187146 63135 187202 63144
rect 187054 59800 187110 59809
rect 187054 59735 187110 59744
rect 186964 53644 187016 53650
rect 186964 53586 187016 53592
rect 186962 49736 187018 49745
rect 186962 49671 187018 49680
rect 186976 41410 187004 49671
rect 187068 45490 187096 59735
rect 187160 48278 187188 63135
rect 187252 60722 187280 86935
rect 187330 83464 187386 83473
rect 187330 83399 187386 83408
rect 187240 60716 187292 60722
rect 187240 60658 187292 60664
rect 187344 57934 187372 83399
rect 187436 82822 187464 130863
rect 188252 130688 188304 130694
rect 188252 130630 188304 130636
rect 188160 130620 188212 130626
rect 188160 130562 188212 130568
rect 187514 124264 187570 124273
rect 187514 124199 187570 124208
rect 187424 82816 187476 82822
rect 187424 82758 187476 82764
rect 187422 80200 187478 80209
rect 187422 80135 187478 80144
rect 187332 57928 187384 57934
rect 187332 57870 187384 57876
rect 187436 56574 187464 80135
rect 187528 80034 187556 124199
rect 187516 80028 187568 80034
rect 187516 79970 187568 79976
rect 187514 76800 187570 76809
rect 187514 76735 187570 76744
rect 187424 56568 187476 56574
rect 187424 56510 187476 56516
rect 187238 56400 187294 56409
rect 187238 56335 187294 56344
rect 187148 48272 187200 48278
rect 187148 48214 187200 48220
rect 187146 46336 187202 46345
rect 187146 46271 187202 46280
rect 187056 45484 187108 45490
rect 187056 45426 187108 45432
rect 186964 41404 187016 41410
rect 186964 41346 187016 41352
rect 186962 39536 187018 39545
rect 186962 39471 187018 39480
rect 186976 35834 187004 39471
rect 187160 38622 187188 46271
rect 187252 44130 187280 56335
rect 187528 55214 187556 76735
rect 187516 55208 187568 55214
rect 187516 55150 187568 55156
rect 187330 53000 187386 53009
rect 187330 52935 187386 52944
rect 187240 44124 187292 44130
rect 187240 44066 187292 44072
rect 187344 42770 187372 52935
rect 187332 42764 187384 42770
rect 187332 42706 187384 42712
rect 187238 40624 187294 40633
rect 187238 40559 187294 40568
rect 187148 38616 187200 38622
rect 187148 38558 187200 38564
rect 187252 35902 187280 40559
rect 187240 35896 187292 35902
rect 187240 35838 187292 35844
rect 186964 35828 187016 35834
rect 186964 35770 187016 35776
rect 186688 30320 186740 30326
rect 186688 30262 186740 30268
rect 182824 28620 182876 28626
rect 182824 28562 182876 28568
rect 188172 28558 188200 130562
rect 188160 28552 188212 28558
rect 188160 28494 188212 28500
rect 188264 28490 188292 130630
rect 188252 28484 188304 28490
rect 188252 28426 188304 28432
rect 188356 28082 188384 297230
rect 188448 29510 188476 297298
rect 188436 29504 188488 29510
rect 188436 29446 188488 29452
rect 188540 29442 188568 297366
rect 190472 267734 190500 304982
rect 190472 267706 190776 267734
rect 190748 249914 190776 267706
rect 193232 249914 193260 306342
rect 204272 267734 204300 325654
rect 207018 307184 207074 307193
rect 207018 307119 207074 307128
rect 207032 306406 207060 307119
rect 207020 306400 207072 306406
rect 207020 306342 207072 306348
rect 207018 305552 207074 305561
rect 207018 305487 207074 305496
rect 207032 305046 207060 305487
rect 207020 305040 207072 305046
rect 207020 304982 207072 304988
rect 204272 267706 204760 267734
rect 201408 256216 201460 256222
rect 201408 256158 201460 256164
rect 195796 253360 195848 253366
rect 195796 253302 195848 253308
rect 195808 249914 195836 253302
rect 198464 253292 198516 253298
rect 198464 253234 198516 253240
rect 198476 249914 198504 253234
rect 201420 252550 201448 256158
rect 202696 254992 202748 254998
rect 202696 254934 202748 254940
rect 200488 252544 200540 252550
rect 200488 252486 200540 252492
rect 201408 252544 201460 252550
rect 201408 252486 201460 252492
rect 200500 249914 200528 252486
rect 190748 249886 191130 249914
rect 193232 249886 193430 249914
rect 195730 249886 195836 249914
rect 198122 249886 198504 249914
rect 200422 249886 200528 249914
rect 202708 249914 202736 254934
rect 204732 249914 204760 267706
rect 207848 254856 207900 254862
rect 207848 254798 207900 254804
rect 207860 249914 207888 254798
rect 208044 253570 208072 327383
rect 208032 253564 208084 253570
rect 208032 253506 208084 253512
rect 208136 253502 208164 328471
rect 208124 253496 208176 253502
rect 208124 253438 208176 253444
rect 208228 253434 208256 329967
rect 208216 253428 208268 253434
rect 208216 253370 208268 253376
rect 208320 253230 208348 334047
rect 209686 332888 209742 332897
rect 209686 332823 209742 332832
rect 209594 331120 209650 331129
rect 209594 331055 209650 331064
rect 209608 254930 209636 331055
rect 209596 254924 209648 254930
rect 209596 254866 209648 254872
rect 209700 254794 209728 332823
rect 238666 299840 238722 299849
rect 238666 299775 238722 299784
rect 215852 298172 215904 298178
rect 215852 298114 215904 298120
rect 215864 298081 215892 298114
rect 215850 298072 215906 298081
rect 215850 298007 215906 298016
rect 224958 298072 225014 298081
rect 224958 298007 225014 298016
rect 226338 298072 226394 298081
rect 226338 298007 226394 298016
rect 227718 298072 227774 298081
rect 227718 298007 227774 298016
rect 229190 298072 229246 298081
rect 229190 298007 229246 298016
rect 230478 298072 230534 298081
rect 230478 298007 230534 298016
rect 231858 298072 231914 298081
rect 231858 298007 231914 298016
rect 233238 298072 233294 298081
rect 233238 298007 233294 298016
rect 234618 298072 234674 298081
rect 234618 298007 234674 298016
rect 237194 298072 237250 298081
rect 237194 298007 237250 298016
rect 219256 256420 219308 256426
rect 219256 256362 219308 256368
rect 210056 256352 210108 256358
rect 210056 256294 210108 256300
rect 209688 254788 209740 254794
rect 209688 254730 209740 254736
rect 208308 253224 208360 253230
rect 208308 253166 208360 253172
rect 210068 249914 210096 256294
rect 212448 256284 212500 256290
rect 212448 256226 212500 256232
rect 212460 249914 212488 256226
rect 217048 255060 217100 255066
rect 217048 255002 217100 255008
rect 214196 253564 214248 253570
rect 214196 253506 214248 253512
rect 202708 249886 202814 249914
rect 204732 249886 205114 249914
rect 207506 249886 207888 249914
rect 209806 249886 210096 249914
rect 212106 249886 212488 249914
rect 214208 249914 214236 253506
rect 217060 249914 217088 255002
rect 219268 249914 219296 256362
rect 221832 253564 221884 253570
rect 221832 253506 221884 253512
rect 221844 249914 221872 253506
rect 223580 253496 223632 253502
rect 223580 253438 223632 253444
rect 214208 249886 214498 249914
rect 216798 249886 217088 249914
rect 219190 249886 219296 249914
rect 221490 249886 221872 249914
rect 223592 249914 223620 253438
rect 224972 253366 225000 298007
rect 226352 256222 226380 298007
rect 227732 297226 227760 298007
rect 227720 297220 227772 297226
rect 227720 297162 227772 297168
rect 227732 256358 227760 297162
rect 229100 297152 229152 297158
rect 229100 297094 229152 297100
rect 227720 256352 227772 256358
rect 227720 256294 227772 256300
rect 226340 256216 226392 256222
rect 226340 256158 226392 256164
rect 229112 253910 229140 297094
rect 229204 297090 229232 298007
rect 229466 297256 229522 297265
rect 229466 297191 229522 297200
rect 229480 297158 229508 297191
rect 229468 297152 229520 297158
rect 229468 297094 229520 297100
rect 229192 297084 229244 297090
rect 229192 297026 229244 297032
rect 229204 256426 229232 297026
rect 229192 256420 229244 256426
rect 229192 256362 229244 256368
rect 230492 254998 230520 298007
rect 231872 256290 231900 298007
rect 231860 256284 231912 256290
rect 231860 256226 231912 256232
rect 230480 254992 230532 254998
rect 230480 254934 230532 254940
rect 228732 253904 228784 253910
rect 228732 253846 228784 253852
rect 229100 253904 229152 253910
rect 229100 253846 229152 253852
rect 226248 253496 226300 253502
rect 226248 253438 226300 253444
rect 224960 253360 225012 253366
rect 224960 253302 225012 253308
rect 226260 249914 226288 253438
rect 228744 249914 228772 253846
rect 233252 253570 233280 298007
rect 233240 253564 233292 253570
rect 233240 253506 233292 253512
rect 232780 253428 232832 253434
rect 232780 253370 232832 253376
rect 231216 253156 231268 253162
rect 231216 253098 231268 253104
rect 231228 249914 231256 253098
rect 223592 249886 223882 249914
rect 226182 249886 226288 249914
rect 228482 249886 228772 249914
rect 230874 249886 231256 249914
rect 232792 249914 232820 253370
rect 234632 253162 234660 298007
rect 237208 253570 237236 298007
rect 237378 297936 237434 297945
rect 237378 297871 237434 297880
rect 237286 297800 237342 297809
rect 237286 297735 237342 297744
rect 237196 253564 237248 253570
rect 237196 253506 237248 253512
rect 235816 253428 235868 253434
rect 235816 253370 235868 253376
rect 234620 253156 234672 253162
rect 234620 253098 234672 253104
rect 235828 249914 235856 253370
rect 237300 252090 237328 297735
rect 237392 253298 237420 297871
rect 238680 297129 238708 299775
rect 243082 299704 243138 299713
rect 243082 299639 243138 299648
rect 238758 298072 238814 298081
rect 238758 298007 238814 298016
rect 240138 298072 240194 298081
rect 240138 298007 240194 298016
rect 241426 298072 241482 298081
rect 241426 298007 241482 298016
rect 242898 298072 242954 298081
rect 242898 298007 242954 298016
rect 238666 297120 238722 297129
rect 238666 297055 238722 297064
rect 238666 296848 238722 296857
rect 238666 296783 238722 296792
rect 237380 253292 237432 253298
rect 237380 253234 237432 253240
rect 238680 252414 238708 296783
rect 238772 254862 238800 298007
rect 240046 297120 240102 297129
rect 240046 297055 240102 297064
rect 238760 254856 238812 254862
rect 238760 254798 238812 254804
rect 240060 253366 240088 297055
rect 240152 255066 240180 298007
rect 240140 255060 240192 255066
rect 240140 255002 240192 255008
rect 240140 254924 240192 254930
rect 240140 254866 240192 254872
rect 240048 253360 240100 253366
rect 240048 253302 240100 253308
rect 238668 252408 238720 252414
rect 238668 252350 238720 252356
rect 237300 252062 237512 252090
rect 232792 249886 233174 249914
rect 235566 249886 235856 249914
rect 237484 249914 237512 252062
rect 240152 249914 240180 254866
rect 241440 252346 241468 298007
rect 241518 297936 241574 297945
rect 241518 297871 241574 297880
rect 241532 253502 241560 297871
rect 242806 297800 242862 297809
rect 242806 297735 242862 297744
rect 242820 256562 242848 297735
rect 242808 256556 242860 256562
rect 242808 256498 242860 256504
rect 242808 253836 242860 253842
rect 242808 253778 242860 253784
rect 241520 253496 241572 253502
rect 241520 253438 241572 253444
rect 241428 252340 241480 252346
rect 241428 252282 241480 252288
rect 242820 249914 242848 253778
rect 242912 253434 242940 298007
rect 243096 297945 243124 299639
rect 244094 298072 244150 298081
rect 244094 298007 244150 298016
rect 244278 298072 244334 298081
rect 244278 298007 244334 298016
rect 245566 298072 245622 298081
rect 245566 298007 245622 298016
rect 246854 298072 246910 298081
rect 246854 298007 246910 298016
rect 248326 298072 248382 298081
rect 248326 298007 248382 298016
rect 249706 298072 249762 298081
rect 249706 298007 249762 298016
rect 251086 298072 251142 298081
rect 251086 298007 251142 298016
rect 252374 298072 252430 298081
rect 252374 298007 252430 298016
rect 253754 298072 253810 298081
rect 253754 298007 253810 298016
rect 255134 298072 255190 298081
rect 255134 298007 255190 298016
rect 256514 298072 256570 298081
rect 256514 298007 256570 298016
rect 257802 298072 257858 298081
rect 257802 298007 257858 298016
rect 257986 298072 258042 298081
rect 257986 298007 258042 298016
rect 259182 298072 259238 298081
rect 259182 298007 259238 298016
rect 260654 298072 260710 298081
rect 260654 298007 260710 298016
rect 262034 298072 262090 298081
rect 262034 298007 262090 298016
rect 263506 298072 263562 298081
rect 263506 298007 263562 298016
rect 266174 298072 266230 298081
rect 266174 298007 266230 298016
rect 273166 298072 273222 298081
rect 273166 298007 273222 298016
rect 274546 298072 274602 298081
rect 274546 298007 274602 298016
rect 275926 298072 275982 298081
rect 275926 298007 275982 298016
rect 277306 298072 277362 298081
rect 277306 298007 277362 298016
rect 243082 297936 243138 297945
rect 243082 297871 243138 297880
rect 244108 254930 244136 298007
rect 244186 297936 244242 297945
rect 244186 297871 244242 297880
rect 244096 254924 244148 254930
rect 244096 254866 244148 254872
rect 242900 253428 242952 253434
rect 242900 253370 242952 253376
rect 244200 253298 244228 297871
rect 244292 253842 244320 298007
rect 245580 257854 245608 298007
rect 246762 297936 246818 297945
rect 246762 297871 246818 297880
rect 246776 259078 246804 297871
rect 246764 259072 246816 259078
rect 246764 259014 246816 259020
rect 245568 257848 245620 257854
rect 245568 257790 245620 257796
rect 244280 253836 244332 253842
rect 244280 253778 244332 253784
rect 246868 253570 246896 298007
rect 248234 297936 248290 297945
rect 248234 297871 248290 297880
rect 246946 297800 247002 297809
rect 246946 297735 247002 297744
rect 246960 253910 246988 297735
rect 248248 259010 248276 297871
rect 248236 259004 248288 259010
rect 248236 258946 248288 258952
rect 247040 254788 247092 254794
rect 247040 254730 247092 254736
rect 246948 253904 247000 253910
rect 246948 253846 247000 253852
rect 244556 253564 244608 253570
rect 244556 253506 244608 253512
rect 246856 253564 246908 253570
rect 246856 253506 246908 253512
rect 244188 253292 244240 253298
rect 244188 253234 244240 253240
rect 237484 249886 237866 249914
rect 240152 249886 240258 249914
rect 242558 249886 242848 249914
rect 244568 249914 244596 253506
rect 247052 249914 247080 254730
rect 248340 253502 248368 298007
rect 249614 297936 249670 297945
rect 249614 297871 249670 297880
rect 249628 258942 249656 297871
rect 249616 258936 249668 258942
rect 249616 258878 249668 258884
rect 249156 253904 249208 253910
rect 249156 253846 249208 253852
rect 248328 253496 248380 253502
rect 248328 253438 248380 253444
rect 249168 249914 249196 253846
rect 249720 253434 249748 298007
rect 250994 297936 251050 297945
rect 250994 297871 251050 297880
rect 251008 258874 251036 297871
rect 250996 258868 251048 258874
rect 250996 258810 251048 258816
rect 250352 256148 250404 256154
rect 250352 256090 250404 256096
rect 249708 253428 249760 253434
rect 249708 253370 249760 253376
rect 250364 252278 250392 256090
rect 251100 254794 251128 298007
rect 252282 297936 252338 297945
rect 252282 297871 252338 297880
rect 252296 258806 252324 297871
rect 252284 258800 252336 258806
rect 252284 258742 252336 258748
rect 252388 254862 252416 298007
rect 252466 297800 252522 297809
rect 252466 297735 252522 297744
rect 252480 255066 252508 297735
rect 253768 260642 253796 298007
rect 253846 297936 253902 297945
rect 253846 297871 253902 297880
rect 253756 260636 253808 260642
rect 253756 260578 253808 260584
rect 252468 255060 252520 255066
rect 252468 255002 252520 255008
rect 253860 254998 253888 297871
rect 255148 260574 255176 298007
rect 255226 297936 255282 297945
rect 255226 297871 255282 297880
rect 255136 260568 255188 260574
rect 255136 260510 255188 260516
rect 255240 256494 255268 297871
rect 256528 260506 256556 298007
rect 256606 297936 256662 297945
rect 256606 297871 256662 297880
rect 256516 260500 256568 260506
rect 256516 260442 256568 260448
rect 255228 256488 255280 256494
rect 255228 256430 255280 256436
rect 256620 256426 256648 297871
rect 257816 260438 257844 298007
rect 257894 297936 257950 297945
rect 257894 297871 257950 297880
rect 257804 260432 257856 260438
rect 257804 260374 257856 260380
rect 256608 256420 256660 256426
rect 256608 256362 256660 256368
rect 257908 256358 257936 297871
rect 257896 256352 257948 256358
rect 257896 256294 257948 256300
rect 258000 256290 258028 298007
rect 259196 261934 259224 298007
rect 259366 297936 259422 297945
rect 259366 297871 259422 297880
rect 259274 297800 259330 297809
rect 259274 297735 259330 297744
rect 259184 261928 259236 261934
rect 259184 261870 259236 261876
rect 259288 260370 259316 297735
rect 259276 260364 259328 260370
rect 259276 260306 259328 260312
rect 257988 256284 258040 256290
rect 257988 256226 258040 256232
rect 259380 256222 259408 297871
rect 260668 260302 260696 298007
rect 260746 297936 260802 297945
rect 260746 297871 260802 297880
rect 260656 260296 260708 260302
rect 260656 260238 260708 260244
rect 260760 257786 260788 297871
rect 262048 258738 262076 298007
rect 262126 297936 262182 297945
rect 262126 297871 262182 297880
rect 263414 297936 263470 297945
rect 263414 297871 263470 297880
rect 262036 258732 262088 258738
rect 262036 258674 262088 258680
rect 260748 257780 260800 257786
rect 260748 257722 260800 257728
rect 262140 257718 262168 297871
rect 263428 261866 263456 297871
rect 263416 261860 263468 261866
rect 263416 261802 263468 261808
rect 262128 257712 262180 257718
rect 262128 257654 262180 257660
rect 263520 257650 263548 298007
rect 264794 296984 264850 296993
rect 264794 296919 264850 296928
rect 264808 261798 264836 296919
rect 264886 296848 264942 296857
rect 264886 296783 264942 296792
rect 264796 261792 264848 261798
rect 264796 261734 264848 261740
rect 263508 257644 263560 257650
rect 263508 257586 263560 257592
rect 259368 256216 259420 256222
rect 259368 256158 259420 256164
rect 253848 254992 253900 254998
rect 253848 254934 253900 254940
rect 252376 254856 252428 254862
rect 252376 254798 252428 254804
rect 251088 254788 251140 254794
rect 251088 254730 251140 254736
rect 264900 253638 264928 296783
rect 266188 261730 266216 298007
rect 269026 297528 269082 297537
rect 269026 297463 269082 297472
rect 267554 297120 267610 297129
rect 267554 297055 267610 297064
rect 266266 296848 266322 296857
rect 266266 296783 266322 296792
rect 267462 296848 267518 296857
rect 267462 296783 267518 296792
rect 266176 261724 266228 261730
rect 266176 261666 266228 261672
rect 266280 257582 266308 296783
rect 267476 263294 267504 296783
rect 267464 263288 267516 263294
rect 267464 263230 267516 263236
rect 267568 261662 267596 297055
rect 267646 296984 267702 296993
rect 267646 296919 267702 296928
rect 267556 261656 267608 261662
rect 267556 261598 267608 261604
rect 266268 257576 266320 257582
rect 266268 257518 266320 257524
rect 264888 253632 264940 253638
rect 264888 253574 264940 253580
rect 267660 253570 267688 296919
rect 268016 256556 268068 256562
rect 268016 256498 268068 256504
rect 256332 253564 256384 253570
rect 256332 253506 256384 253512
rect 267648 253564 267700 253570
rect 267648 253506 267700 253512
rect 253940 253224 253992 253230
rect 253940 253166 253992 253172
rect 251548 252408 251600 252414
rect 251548 252350 251600 252356
rect 250352 252272 250404 252278
rect 250352 252214 250404 252220
rect 251560 249914 251588 252350
rect 253952 249914 253980 253166
rect 256344 249914 256372 253506
rect 260932 253496 260984 253502
rect 260932 253438 260984 253444
rect 258540 253360 258592 253366
rect 258540 253302 258592 253308
rect 258552 249914 258580 253302
rect 260944 249914 260972 253438
rect 265532 253428 265584 253434
rect 265532 253370 265584 253376
rect 263692 252340 263744 252346
rect 263692 252282 263744 252288
rect 263704 249914 263732 252282
rect 244568 249886 244950 249914
rect 247052 249886 247250 249914
rect 249168 249886 249550 249914
rect 251560 249886 251942 249914
rect 253952 249886 254242 249914
rect 256344 249886 256634 249914
rect 258552 249886 258934 249914
rect 260944 249886 261326 249914
rect 263626 249886 263732 249914
rect 265544 249914 265572 253370
rect 268028 249914 268056 256498
rect 269040 253502 269068 297463
rect 270406 296848 270462 296857
rect 270406 296783 270462 296792
rect 271786 296848 271842 296857
rect 271786 296783 271842 296792
rect 273074 296848 273130 296857
rect 273074 296783 273130 296792
rect 269028 253496 269080 253502
rect 269028 253438 269080 253444
rect 270420 253434 270448 296783
rect 270500 254788 270552 254794
rect 270500 254730 270552 254736
rect 270408 253428 270460 253434
rect 270408 253370 270460 253376
rect 270512 249914 270540 254730
rect 271800 253366 271828 296783
rect 273088 257514 273116 296783
rect 273076 257508 273128 257514
rect 273076 257450 273128 257456
rect 273180 254794 273208 298007
rect 273168 254788 273220 254794
rect 273168 254730 273220 254736
rect 271788 253360 271840 253366
rect 271788 253302 271840 253308
rect 274560 253298 274588 298007
rect 274916 255060 274968 255066
rect 274916 255002 274968 255008
rect 272708 253292 272760 253298
rect 272708 253234 272760 253240
rect 274548 253292 274600 253298
rect 274548 253234 274600 253240
rect 272720 249914 272748 253234
rect 274928 249914 274956 255002
rect 275940 253230 275968 298007
rect 277320 256154 277348 298007
rect 352564 297016 352616 297022
rect 352564 296958 352616 296964
rect 338120 261928 338172 261934
rect 338120 261870 338172 261876
rect 314752 260636 314804 260642
rect 314752 260578 314804 260584
rect 286600 259072 286652 259078
rect 286600 259014 286652 259020
rect 282092 257848 282144 257854
rect 282092 257790 282144 257796
rect 277308 256148 277360 256154
rect 277308 256090 277360 256096
rect 279700 254992 279752 254998
rect 279700 254934 279752 254940
rect 277492 254924 277544 254930
rect 277492 254866 277544 254872
rect 275928 253224 275980 253230
rect 275928 253166 275980 253172
rect 277504 249914 277532 254866
rect 279712 249914 279740 254934
rect 282104 249914 282132 257790
rect 284300 256488 284352 256494
rect 284300 256430 284352 256436
rect 284312 249914 284340 256430
rect 286612 249914 286640 259014
rect 291200 259004 291252 259010
rect 291200 258946 291252 258952
rect 289084 256420 289136 256426
rect 289084 256362 289136 256368
rect 289096 249914 289124 256362
rect 291212 249914 291240 258946
rect 295984 258936 296036 258942
rect 295984 258878 296036 258884
rect 293960 256352 294012 256358
rect 293960 256294 294012 256300
rect 293972 249914 294000 256294
rect 295996 249914 296024 258878
rect 300860 258868 300912 258874
rect 300860 258810 300912 258816
rect 298468 256284 298520 256290
rect 298468 256226 298520 256232
rect 298480 249914 298508 256226
rect 300872 249914 300900 258810
rect 305368 258800 305420 258806
rect 305368 258742 305420 258748
rect 303068 256216 303120 256222
rect 303068 256158 303120 256164
rect 303080 249914 303108 256158
rect 305380 249914 305408 258742
rect 307760 257780 307812 257786
rect 307760 257722 307812 257728
rect 307772 249914 307800 257722
rect 312452 257712 312504 257718
rect 312452 257654 312504 257660
rect 310060 254856 310112 254862
rect 310060 254798 310112 254804
rect 310072 249914 310100 254798
rect 312464 249914 312492 257654
rect 314764 249914 314792 260578
rect 319352 260568 319404 260574
rect 319352 260510 319404 260516
rect 317512 257644 317564 257650
rect 317512 257586 317564 257592
rect 317524 249914 317552 257586
rect 265544 249886 265926 249914
rect 268028 249886 268318 249914
rect 270512 249886 270618 249914
rect 272720 249886 273010 249914
rect 274928 249886 275310 249914
rect 277504 249886 277702 249914
rect 279712 249886 280002 249914
rect 282104 249886 282394 249914
rect 284312 249886 284694 249914
rect 286612 249886 286994 249914
rect 289096 249886 289386 249914
rect 291212 249886 291686 249914
rect 293972 249886 294078 249914
rect 295996 249886 296378 249914
rect 298480 249886 298770 249914
rect 300872 249886 301070 249914
rect 303080 249886 303370 249914
rect 305380 249886 305762 249914
rect 307772 249886 308062 249914
rect 310072 249886 310454 249914
rect 312464 249886 312754 249914
rect 314764 249886 315146 249914
rect 317446 249886 317552 249914
rect 319364 249914 319392 260510
rect 324320 260500 324372 260506
rect 324320 260442 324372 260448
rect 321836 253632 321888 253638
rect 321836 253574 321888 253580
rect 321848 249914 321876 253574
rect 324332 249914 324360 260442
rect 328736 260432 328788 260438
rect 328736 260374 328788 260380
rect 326436 257576 326488 257582
rect 326436 257518 326488 257524
rect 326448 249914 326476 257518
rect 328748 249914 328776 260374
rect 333336 260364 333388 260370
rect 333336 260306 333388 260312
rect 331220 253564 331272 253570
rect 331220 253506 331272 253512
rect 331232 249914 331260 253506
rect 333348 249914 333376 260306
rect 335820 253496 335872 253502
rect 335820 253438 335872 253444
rect 335832 249914 335860 253438
rect 338132 249914 338160 261870
rect 352104 261860 352156 261866
rect 352104 261802 352156 261808
rect 342720 260296 342772 260302
rect 342720 260238 342772 260244
rect 340420 253428 340472 253434
rect 340420 253370 340472 253376
rect 340432 249914 340460 253370
rect 342732 249914 342760 260238
rect 347780 258732 347832 258738
rect 347780 258674 347832 258680
rect 345204 253360 345256 253366
rect 345204 253302 345256 253308
rect 345216 249914 345244 253302
rect 347792 249914 347820 258674
rect 349804 254788 349856 254794
rect 349804 254730 349856 254736
rect 349816 249914 349844 254730
rect 352116 249914 352144 261802
rect 352576 252346 352604 296958
rect 409144 296948 409196 296954
rect 409144 296890 409196 296896
rect 409052 296880 409104 296886
rect 409052 296822 409104 296828
rect 408960 296812 409012 296818
rect 408960 296754 409012 296760
rect 408868 296744 408920 296750
rect 408868 296686 408920 296692
rect 371332 263288 371384 263294
rect 371332 263230 371384 263236
rect 356704 261792 356756 261798
rect 356704 261734 356756 261740
rect 354772 257508 354824 257514
rect 354772 257450 354824 257456
rect 352564 252340 352616 252346
rect 352564 252282 352616 252288
rect 354784 249914 354812 257450
rect 356716 249914 356744 261734
rect 361580 261724 361632 261730
rect 361580 261666 361632 261672
rect 359188 253292 359240 253298
rect 359188 253234 359240 253240
rect 359200 249914 359228 253234
rect 361592 249914 361620 261666
rect 366088 261656 366140 261662
rect 366088 261598 366140 261604
rect 363972 253224 364024 253230
rect 363972 253166 364024 253172
rect 363984 249914 364012 253166
rect 366100 249914 366128 261598
rect 368572 256148 368624 256154
rect 368572 256090 368624 256096
rect 368584 249914 368612 256090
rect 371344 249914 371372 263230
rect 406016 261588 406068 261594
rect 406016 261530 406068 261536
rect 385040 261520 385092 261526
rect 385040 261462 385092 261468
rect 378140 260228 378192 260234
rect 378140 260170 378192 260176
rect 373356 254720 373408 254726
rect 373356 254662 373408 254668
rect 319364 249886 319746 249914
rect 321848 249886 322138 249914
rect 324332 249886 324438 249914
rect 326448 249886 326830 249914
rect 328748 249886 329130 249914
rect 331232 249886 331522 249914
rect 333348 249886 333822 249914
rect 335832 249886 336214 249914
rect 338132 249886 338514 249914
rect 340432 249886 340814 249914
rect 342732 249886 343206 249914
rect 345216 249886 345506 249914
rect 347792 249886 347898 249914
rect 349816 249886 350198 249914
rect 352116 249886 352590 249914
rect 354784 249886 354890 249914
rect 356716 249886 357190 249914
rect 359200 249886 359582 249914
rect 361592 249886 361882 249914
rect 363984 249886 364274 249914
rect 366100 249886 366574 249914
rect 368584 249886 368966 249914
rect 371266 249886 371372 249914
rect 373368 249914 373396 254662
rect 375564 251864 375616 251870
rect 375564 251806 375616 251812
rect 375576 249914 375604 251806
rect 378152 249914 378180 260170
rect 382556 254652 382608 254658
rect 382556 254594 382608 254600
rect 382568 249914 382596 254594
rect 385052 249914 385080 261462
rect 401600 260160 401652 260166
rect 401600 260102 401652 260108
rect 387340 256080 387392 256086
rect 387340 256022 387392 256028
rect 387352 249914 387380 256022
rect 394332 252340 394384 252346
rect 394332 252282 394384 252288
rect 391940 252204 391992 252210
rect 391940 252146 391992 252152
rect 389732 252068 389784 252074
rect 389732 252010 389784 252016
rect 389744 249914 389772 252010
rect 391952 249914 391980 252146
rect 394344 249914 394372 252282
rect 398932 252000 398984 252006
rect 398932 251942 398984 251948
rect 396724 251932 396776 251938
rect 396724 251874 396776 251880
rect 396736 249914 396764 251874
rect 398944 249914 398972 251942
rect 401612 249914 401640 260102
rect 403716 252272 403768 252278
rect 403716 252214 403768 252220
rect 403728 249914 403756 252214
rect 406028 249914 406056 261530
rect 408592 252136 408644 252142
rect 408592 252078 408644 252084
rect 408500 250844 408552 250850
rect 408500 250786 408552 250792
rect 373368 249886 373658 249914
rect 375576 249886 375958 249914
rect 378152 249886 378258 249914
rect 382568 249886 382950 249914
rect 385052 249886 385342 249914
rect 387352 249886 387642 249914
rect 389744 249886 390034 249914
rect 391952 249886 392334 249914
rect 394344 249886 394634 249914
rect 396736 249886 397026 249914
rect 398944 249886 399326 249914
rect 401612 249886 401718 249914
rect 403728 249886 404018 249914
rect 406028 249886 406410 249914
rect 408512 249665 408540 250786
rect 408604 249914 408632 252078
rect 408604 249886 408710 249914
rect 408498 249656 408554 249665
rect 408498 249591 408554 249600
rect 408880 230058 408908 296686
rect 408972 231826 409000 296754
rect 409064 238754 409092 296822
rect 409156 267734 409184 296890
rect 409156 267706 409368 267734
rect 409340 247761 409368 267706
rect 411628 263220 411680 263226
rect 411628 263162 411680 263168
rect 410432 263152 410484 263158
rect 410432 263094 410484 263100
rect 409972 263016 410024 263022
rect 409972 262958 410024 262964
rect 409880 257372 409932 257378
rect 409880 257314 409932 257320
rect 409326 247752 409382 247761
rect 409326 247687 409382 247696
rect 409064 238726 409368 238754
rect 409340 233753 409368 238726
rect 409326 233744 409382 233753
rect 409326 233679 409382 233688
rect 409326 231840 409382 231849
rect 408972 231798 409326 231826
rect 409326 231775 409382 231784
rect 409326 230072 409382 230081
rect 408880 230030 409326 230058
rect 409326 230007 409382 230016
rect 409892 212401 409920 257314
rect 409984 223281 410012 262958
rect 410064 262948 410116 262954
rect 410064 262890 410116 262896
rect 410076 226137 410104 262890
rect 410340 257440 410392 257446
rect 410340 257382 410392 257388
rect 410248 256012 410300 256018
rect 410248 255954 410300 255960
rect 410156 254584 410208 254590
rect 410156 254526 410208 254532
rect 410062 226128 410118 226137
rect 410062 226063 410118 226072
rect 409970 223272 410026 223281
rect 409970 223207 410026 223216
rect 410168 217705 410196 254526
rect 410260 221649 410288 255954
rect 410352 227497 410380 257382
rect 410444 241233 410472 263094
rect 411536 263084 411588 263090
rect 411536 263026 411588 263032
rect 410524 250776 410576 250782
rect 410524 250718 410576 250724
rect 410536 243273 410564 250718
rect 411260 250708 411312 250714
rect 411260 250650 411312 250656
rect 411272 245177 411300 250650
rect 411444 250640 411496 250646
rect 411444 250582 411496 250588
rect 411352 250504 411404 250510
rect 411352 250446 411404 250452
rect 411258 245168 411314 245177
rect 411258 245103 411314 245112
rect 411260 243568 411312 243574
rect 411260 243510 411312 243516
rect 410522 243264 410578 243273
rect 410522 243199 410578 243208
rect 410430 241224 410486 241233
rect 410430 241159 410486 241168
rect 411272 235385 411300 243510
rect 411258 235376 411314 235385
rect 411258 235311 411314 235320
rect 410338 227488 410394 227497
rect 410338 227423 410394 227432
rect 410246 221640 410302 221649
rect 410246 221575 410302 221584
rect 410154 217696 410210 217705
rect 410154 217631 410210 217640
rect 411364 213761 411392 250446
rect 411456 243574 411484 250582
rect 411444 243568 411496 243574
rect 411444 243510 411496 243516
rect 411444 243432 411496 243438
rect 411444 243374 411496 243380
rect 411456 215665 411484 243374
rect 411548 237289 411576 263026
rect 411640 239329 411668 263162
rect 411720 262880 411772 262886
rect 411720 262822 411772 262828
rect 411626 239320 411682 239329
rect 411626 239255 411682 239264
rect 411534 237280 411590 237289
rect 411534 237215 411590 237224
rect 411732 219609 411760 262822
rect 411812 250572 411864 250578
rect 411812 250514 411864 250520
rect 411824 243438 411852 250514
rect 580356 249824 580408 249830
rect 580356 249766 580408 249772
rect 580264 248464 580316 248470
rect 580264 248406 580316 248412
rect 411812 243432 411864 243438
rect 411812 243374 411864 243380
rect 579618 232384 579674 232393
rect 579618 232319 579674 232328
rect 579632 231878 579660 232319
rect 463700 231872 463752 231878
rect 463700 231814 463752 231820
rect 579620 231872 579672 231878
rect 579620 231814 579672 231820
rect 411718 219600 411774 219609
rect 411718 219535 411774 219544
rect 411442 215656 411498 215665
rect 411442 215591 411498 215600
rect 411350 213752 411406 213761
rect 411350 213687 411406 213696
rect 409878 212392 409934 212401
rect 409878 212327 409934 212336
rect 411260 209840 411312 209846
rect 411258 209808 411260 209817
rect 418804 209840 418856 209846
rect 411312 209808 411314 209817
rect 418804 209782 418856 209788
rect 411258 209743 411314 209752
rect 411258 207904 411314 207913
rect 411258 207839 411314 207848
rect 411272 207058 411300 207839
rect 411260 207052 411312 207058
rect 411260 206994 411312 207000
rect 414664 207052 414716 207058
rect 414664 206994 414716 207000
rect 411258 205864 411314 205873
rect 411258 205799 411314 205808
rect 411272 205698 411300 205799
rect 411260 205692 411312 205698
rect 411260 205634 411312 205640
rect 411258 203960 411314 203969
rect 411258 203895 411314 203904
rect 411272 202910 411300 203895
rect 411260 202904 411312 202910
rect 411260 202846 411312 202852
rect 411902 201920 411958 201929
rect 411902 201855 411958 201864
rect 411258 197976 411314 197985
rect 411258 197911 411314 197920
rect 411272 197402 411300 197911
rect 411260 197396 411312 197402
rect 411260 197338 411312 197344
rect 411258 196072 411314 196081
rect 411258 196007 411260 196016
rect 411312 196007 411314 196016
rect 411260 195978 411312 195984
rect 411258 192128 411314 192137
rect 411258 192063 411314 192072
rect 411272 191894 411300 192063
rect 411260 191888 411312 191894
rect 411260 191830 411312 191836
rect 411258 190224 411314 190233
rect 411258 190159 411314 190168
rect 411272 189106 411300 190159
rect 411260 189100 411312 189106
rect 411260 189042 411312 189048
rect 411258 188184 411314 188193
rect 411258 188119 411314 188128
rect 411272 187746 411300 188119
rect 411260 187740 411312 187746
rect 411260 187682 411312 187688
rect 411258 186280 411314 186289
rect 411258 186215 411314 186224
rect 411272 184958 411300 186215
rect 411260 184952 411312 184958
rect 411260 184894 411312 184900
rect 411258 184240 411314 184249
rect 411258 184175 411314 184184
rect 411272 183598 411300 184175
rect 411260 183592 411312 183598
rect 411260 183534 411312 183540
rect 411258 182336 411314 182345
rect 411258 182271 411314 182280
rect 411272 182238 411300 182271
rect 411260 182232 411312 182238
rect 411260 182174 411312 182180
rect 411258 180296 411314 180305
rect 411258 180231 411314 180240
rect 411272 179450 411300 180231
rect 411260 179444 411312 179450
rect 411260 179386 411312 179392
rect 411258 178392 411314 178401
rect 411258 178327 411314 178336
rect 411272 178090 411300 178327
rect 411260 178084 411312 178090
rect 411260 178026 411312 178032
rect 411258 176488 411314 176497
rect 411258 176423 411314 176432
rect 411272 175302 411300 176423
rect 411260 175296 411312 175302
rect 411260 175238 411312 175244
rect 411258 174448 411314 174457
rect 411258 174383 411314 174392
rect 411272 173942 411300 174383
rect 411260 173936 411312 173942
rect 411260 173878 411312 173884
rect 411260 172576 411312 172582
rect 411258 172544 411260 172553
rect 411312 172544 411314 172553
rect 411258 172479 411314 172488
rect 411258 170504 411314 170513
rect 411258 170439 411314 170448
rect 411272 169794 411300 170439
rect 411260 169788 411312 169794
rect 411260 169730 411312 169736
rect 411258 168600 411314 168609
rect 411258 168535 411314 168544
rect 411272 168434 411300 168535
rect 411260 168428 411312 168434
rect 411260 168370 411312 168376
rect 411258 166560 411314 166569
rect 411258 166495 411314 166504
rect 411272 165646 411300 166495
rect 411260 165640 411312 165646
rect 411260 165582 411312 165588
rect 411258 164656 411314 164665
rect 411258 164591 411314 164600
rect 411272 164286 411300 164591
rect 411260 164280 411312 164286
rect 411260 164222 411312 164228
rect 411258 162616 411314 162625
rect 411258 162551 411314 162560
rect 411272 161498 411300 162551
rect 411260 161492 411312 161498
rect 411260 161434 411312 161440
rect 411258 160712 411314 160721
rect 411258 160647 411314 160656
rect 411272 160138 411300 160647
rect 411260 160132 411312 160138
rect 411260 160074 411312 160080
rect 411258 158808 411314 158817
rect 411258 158743 411260 158752
rect 411312 158743 411314 158752
rect 411260 158714 411312 158720
rect 411258 156768 411314 156777
rect 411258 156703 411314 156712
rect 411272 155990 411300 156703
rect 411260 155984 411312 155990
rect 411260 155926 411312 155932
rect 411258 154864 411314 154873
rect 411258 154799 411314 154808
rect 411272 154630 411300 154799
rect 411260 154624 411312 154630
rect 411260 154566 411312 154572
rect 411258 152824 411314 152833
rect 411258 152759 411314 152768
rect 411272 151842 411300 152759
rect 411260 151836 411312 151842
rect 411260 151778 411312 151784
rect 411258 150920 411314 150929
rect 411258 150855 411314 150864
rect 411272 150482 411300 150855
rect 411260 150476 411312 150482
rect 411260 150418 411312 150424
rect 411258 148880 411314 148889
rect 411258 148815 411314 148824
rect 411272 147694 411300 148815
rect 411260 147688 411312 147694
rect 411260 147630 411312 147636
rect 411258 146976 411314 146985
rect 411258 146911 411314 146920
rect 411272 146334 411300 146911
rect 411260 146328 411312 146334
rect 411260 146270 411312 146276
rect 411260 144968 411312 144974
rect 411258 144936 411260 144945
rect 411312 144936 411314 144945
rect 411258 144871 411314 144880
rect 411258 143032 411314 143041
rect 411258 142967 411314 142976
rect 411272 142186 411300 142967
rect 411260 142180 411312 142186
rect 411260 142122 411312 142128
rect 411258 141128 411314 141137
rect 411258 141063 411314 141072
rect 411272 140826 411300 141063
rect 411260 140820 411312 140826
rect 411260 140762 411312 140768
rect 411258 139088 411314 139097
rect 411258 139023 411314 139032
rect 411272 138038 411300 139023
rect 411260 138032 411312 138038
rect 411260 137974 411312 137980
rect 411258 137184 411314 137193
rect 411258 137119 411314 137128
rect 411272 136678 411300 137119
rect 411260 136672 411312 136678
rect 411260 136614 411312 136620
rect 411258 135144 411314 135153
rect 411258 135079 411314 135088
rect 411272 133958 411300 135079
rect 411260 133952 411312 133958
rect 411260 133894 411312 133900
rect 411258 133240 411314 133249
rect 411258 133175 411314 133184
rect 411272 132530 411300 133175
rect 411260 132524 411312 132530
rect 411260 132466 411312 132472
rect 188712 132116 188764 132122
rect 188712 132058 188764 132064
rect 188620 131776 188672 131782
rect 188620 131718 188672 131724
rect 188528 29436 188580 29442
rect 188528 29378 188580 29384
rect 188632 28286 188660 131718
rect 188724 28830 188752 132058
rect 188988 132048 189040 132054
rect 188988 131990 189040 131996
rect 188804 131912 188856 131918
rect 188804 131854 188856 131860
rect 188712 28824 188764 28830
rect 188712 28766 188764 28772
rect 188816 28422 188844 131854
rect 188896 131844 188948 131850
rect 188896 131786 188948 131792
rect 188908 28762 188936 131786
rect 188896 28756 188948 28762
rect 188896 28698 188948 28704
rect 189000 28694 189028 131990
rect 410524 131436 410576 131442
rect 410524 131378 410576 131384
rect 189816 130552 189868 130558
rect 189868 130500 189948 130506
rect 189816 130494 189948 130500
rect 189724 130484 189776 130490
rect 189828 130478 189948 130494
rect 189724 130426 189776 130432
rect 188988 28688 189040 28694
rect 188988 28630 189040 28636
rect 188804 28416 188856 28422
rect 188804 28358 188856 28364
rect 188620 28280 188672 28286
rect 188620 28222 188672 28228
rect 189736 28150 189764 130426
rect 189816 130416 189868 130422
rect 189816 130358 189868 130364
rect 189828 28354 189856 130358
rect 189816 28348 189868 28354
rect 189816 28290 189868 28296
rect 189920 28218 189948 130478
rect 194074 30110 194456 30138
rect 202170 30110 202552 30138
rect 210358 30110 210648 30138
rect 194428 29238 194456 30110
rect 202524 29306 202552 30110
rect 201500 29300 201552 29306
rect 201500 29242 201552 29248
rect 202512 29300 202564 29306
rect 202512 29242 202564 29248
rect 193220 29232 193272 29238
rect 193220 29174 193272 29180
rect 194416 29232 194468 29238
rect 194416 29174 194468 29180
rect 189908 28212 189960 28218
rect 189908 28154 189960 28160
rect 189724 28144 189776 28150
rect 189724 28086 189776 28092
rect 188344 28076 188396 28082
rect 188344 28018 188396 28024
rect 79968 27600 80020 27606
rect 79968 27542 80020 27548
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 1308 4072 1360 4078
rect 1308 4014 1360 4020
rect 1320 3670 1348 4014
rect 2700 3738 2728 4082
rect 193232 4078 193260 29174
rect 201512 4146 201540 29242
rect 210620 29034 210648 30110
rect 218072 30110 218454 30138
rect 226642 30110 227024 30138
rect 210608 29028 210660 29034
rect 210608 28970 210660 28976
rect 218072 6866 218100 30110
rect 226996 29102 227024 30110
rect 234632 30110 234738 30138
rect 242926 30110 243032 30138
rect 226984 29096 227036 29102
rect 226984 29038 227036 29044
rect 234632 28082 234660 30110
rect 243004 29374 243032 30110
rect 258920 30110 259210 30138
rect 267016 30110 267398 30138
rect 275112 30110 275494 30138
rect 283392 30110 283682 30138
rect 299584 30110 299966 30138
rect 307772 30110 308062 30138
rect 316144 30110 316250 30138
rect 324346 30110 324452 30138
rect 258920 29510 258948 30110
rect 258908 29504 258960 29510
rect 258908 29446 258960 29452
rect 242992 29368 243044 29374
rect 242992 29310 243044 29316
rect 267016 28150 267044 30110
rect 275112 28218 275140 30110
rect 283392 28286 283420 30110
rect 299584 29442 299612 30110
rect 299572 29436 299624 29442
rect 299572 29378 299624 29384
rect 307772 28354 307800 30110
rect 316144 28422 316172 30110
rect 324424 28490 324452 30110
rect 332152 30110 332534 30138
rect 340432 30110 340722 30138
rect 348528 30110 348818 30138
rect 356624 30110 357006 30138
rect 364720 30110 365102 30138
rect 373000 30110 373290 30138
rect 381096 30110 381386 30138
rect 389192 30110 389574 30138
rect 397472 30110 397670 30138
rect 405752 30110 405858 30138
rect 332152 28558 332180 30110
rect 340432 28626 340460 30110
rect 348528 28694 348556 30110
rect 356624 28762 356652 30110
rect 364720 29170 364748 30110
rect 364708 29164 364760 29170
rect 364708 29106 364760 29112
rect 373000 28898 373028 30110
rect 381096 28966 381124 30110
rect 381084 28960 381136 28966
rect 381084 28902 381136 28908
rect 372988 28892 373040 28898
rect 372988 28834 373040 28840
rect 389192 28830 389220 30110
rect 389180 28824 389232 28830
rect 397472 28801 397500 30110
rect 405752 28937 405780 30110
rect 410536 29238 410564 131378
rect 411258 129296 411314 129305
rect 411258 129231 411314 129240
rect 411272 128518 411300 129231
rect 411260 128512 411312 128518
rect 411260 128454 411312 128460
rect 411258 127256 411314 127265
rect 411258 127191 411314 127200
rect 411272 127090 411300 127191
rect 411260 127084 411312 127090
rect 411260 127026 411312 127032
rect 411258 125352 411314 125361
rect 411258 125287 411314 125296
rect 411272 124302 411300 125287
rect 411260 124296 411312 124302
rect 411260 124238 411312 124244
rect 411258 123312 411314 123321
rect 411258 123247 411314 123256
rect 411272 122942 411300 123247
rect 411260 122936 411312 122942
rect 411260 122878 411312 122884
rect 411258 121408 411314 121417
rect 411258 121343 411314 121352
rect 410616 120760 410668 120766
rect 410616 120702 410668 120708
rect 410628 29306 410656 120702
rect 411272 120154 411300 121343
rect 411260 120148 411312 120154
rect 411260 120090 411312 120096
rect 411258 119504 411314 119513
rect 411258 119439 411314 119448
rect 411272 118726 411300 119439
rect 411260 118720 411312 118726
rect 411260 118662 411312 118668
rect 411258 115560 411314 115569
rect 411258 115495 411314 115504
rect 411272 114578 411300 115495
rect 411260 114572 411312 114578
rect 411260 114514 411312 114520
rect 411916 114510 411944 201855
rect 412086 200016 412142 200025
rect 412086 199951 412142 199960
rect 411994 194168 412050 194177
rect 411994 194103 412050 194112
rect 411904 114504 411956 114510
rect 411904 114446 411956 114452
rect 411258 113520 411314 113529
rect 411258 113455 411314 113464
rect 411272 113218 411300 113455
rect 411260 113212 411312 113218
rect 411260 113154 411312 113160
rect 411902 111616 411958 111625
rect 411902 111551 411958 111560
rect 411258 109576 411314 109585
rect 411258 109511 411314 109520
rect 411272 109070 411300 109511
rect 411260 109064 411312 109070
rect 411260 109006 411312 109012
rect 411260 107704 411312 107710
rect 411258 107672 411260 107681
rect 411312 107672 411314 107681
rect 411258 107607 411314 107616
rect 411258 103728 411314 103737
rect 411258 103663 411314 103672
rect 411272 103562 411300 103663
rect 411260 103556 411312 103562
rect 411260 103498 411312 103504
rect 411258 101824 411314 101833
rect 411258 101759 411314 101768
rect 411272 100774 411300 101759
rect 411260 100768 411312 100774
rect 411260 100710 411312 100716
rect 411260 95872 411312 95878
rect 411258 95840 411260 95849
rect 411312 95840 411314 95849
rect 411258 95775 411314 95784
rect 411260 93968 411312 93974
rect 411258 93936 411260 93945
rect 411312 93936 411314 93945
rect 411258 93871 411314 93880
rect 411260 92472 411312 92478
rect 411260 92414 411312 92420
rect 411272 91905 411300 92414
rect 411258 91896 411314 91905
rect 411258 91831 411314 91840
rect 411258 89992 411314 90001
rect 411258 89927 411314 89936
rect 411272 89826 411300 89927
rect 411260 89820 411312 89826
rect 411260 89762 411312 89768
rect 411260 88324 411312 88330
rect 411260 88266 411312 88272
rect 411272 87961 411300 88266
rect 411258 87952 411314 87961
rect 411258 87887 411314 87896
rect 411260 86488 411312 86494
rect 411260 86430 411312 86436
rect 411272 86057 411300 86430
rect 411258 86048 411314 86057
rect 411258 85983 411314 85992
rect 411260 84176 411312 84182
rect 411258 84144 411260 84153
rect 411312 84144 411314 84153
rect 411258 84079 411314 84088
rect 411258 82104 411314 82113
rect 411258 82039 411314 82048
rect 411272 81462 411300 82039
rect 411260 81456 411312 81462
rect 411260 81398 411312 81404
rect 411260 78260 411312 78266
rect 411260 78202 411312 78208
rect 411272 78169 411300 78202
rect 411258 78160 411314 78169
rect 411258 78095 411314 78104
rect 411260 76764 411312 76770
rect 411260 76706 411312 76712
rect 411272 76265 411300 76706
rect 411258 76256 411314 76265
rect 411258 76191 411314 76200
rect 411260 74248 411312 74254
rect 411258 74216 411260 74225
rect 411312 74216 411314 74225
rect 411258 74151 411314 74160
rect 411260 73160 411312 73166
rect 411260 73102 411312 73108
rect 411272 72321 411300 73102
rect 411258 72312 411314 72321
rect 411258 72247 411314 72256
rect 411350 70272 411406 70281
rect 411350 70207 411406 70216
rect 411364 69086 411392 70207
rect 411352 69080 411404 69086
rect 411352 69022 411404 69028
rect 411260 69012 411312 69018
rect 411260 68954 411312 68960
rect 411272 68377 411300 68954
rect 411258 68368 411314 68377
rect 411258 68303 411314 68312
rect 411258 66464 411314 66473
rect 411258 66399 411314 66408
rect 411272 66298 411300 66399
rect 411260 66292 411312 66298
rect 411260 66234 411312 66240
rect 411260 64524 411312 64530
rect 411260 64466 411312 64472
rect 411272 64433 411300 64466
rect 411258 64424 411314 64433
rect 411258 64359 411314 64368
rect 411260 63504 411312 63510
rect 411260 63446 411312 63452
rect 411272 62529 411300 63446
rect 411258 62520 411314 62529
rect 411258 62455 411314 62464
rect 411258 60480 411314 60489
rect 411258 60415 411314 60424
rect 411272 59430 411300 60415
rect 411260 59424 411312 59430
rect 411260 59366 411312 59372
rect 411258 58576 411314 58585
rect 411258 58511 411314 58520
rect 411272 58002 411300 58511
rect 411260 57996 411312 58002
rect 411260 57938 411312 57944
rect 411258 54632 411314 54641
rect 411258 54567 411314 54576
rect 411272 54058 411300 54567
rect 411260 54052 411312 54058
rect 411260 53994 411312 54000
rect 411258 52592 411314 52601
rect 411258 52527 411260 52536
rect 411312 52527 411314 52536
rect 411260 52498 411312 52504
rect 411258 48784 411314 48793
rect 411258 48719 411314 48728
rect 411272 48346 411300 48719
rect 411260 48340 411312 48346
rect 411260 48282 411312 48288
rect 411258 42800 411314 42809
rect 411916 42770 411944 111551
rect 412008 107642 412036 194103
rect 412100 113150 412128 199951
rect 414676 139398 414704 206994
rect 416044 196036 416096 196042
rect 416044 195978 416096 195984
rect 414940 151836 414992 151842
rect 414940 151778 414992 151784
rect 414664 139392 414716 139398
rect 414664 139334 414716 139340
rect 414664 131368 414716 131374
rect 414664 131310 414716 131316
rect 412178 131200 412234 131209
rect 412178 131135 412234 131144
rect 412088 113144 412140 113150
rect 412088 113086 412140 113092
rect 411996 107636 412048 107642
rect 411996 107578 412048 107584
rect 411994 105632 412050 105641
rect 411994 105567 412050 105576
rect 411258 42735 411314 42744
rect 411904 42764 411956 42770
rect 411272 42702 411300 42735
rect 411904 42706 411956 42712
rect 411260 42696 411312 42702
rect 411260 42638 411312 42644
rect 411260 41064 411312 41070
rect 411260 41006 411312 41012
rect 411272 40905 411300 41006
rect 411258 40896 411314 40905
rect 411258 40831 411314 40840
rect 411904 40724 411956 40730
rect 411904 40666 411956 40672
rect 411260 38888 411312 38894
rect 411258 38856 411260 38865
rect 411312 38856 411314 38865
rect 411258 38791 411314 38800
rect 411260 37188 411312 37194
rect 411260 37130 411312 37136
rect 411272 36961 411300 37130
rect 411258 36952 411314 36961
rect 411258 36887 411314 36896
rect 411260 35828 411312 35834
rect 411260 35770 411312 35776
rect 411272 34921 411300 35770
rect 411258 34912 411314 34921
rect 411258 34847 411314 34856
rect 411260 33108 411312 33114
rect 411260 33050 411312 33056
rect 411272 33017 411300 33050
rect 411258 33008 411314 33017
rect 411258 32943 411314 32952
rect 411258 31104 411314 31113
rect 411258 31039 411314 31048
rect 411272 30258 411300 31039
rect 411260 30252 411312 30258
rect 411260 30194 411312 30200
rect 411916 30190 411944 40666
rect 412008 37262 412036 105567
rect 412086 99784 412142 99793
rect 412086 99719 412142 99728
rect 411996 37256 412048 37262
rect 411996 37198 412048 37204
rect 412100 33046 412128 99719
rect 412192 57934 412220 131135
rect 413284 130008 413336 130014
rect 413284 129950 413336 129956
rect 412456 128376 412508 128382
rect 412456 128318 412508 128324
rect 412270 117464 412326 117473
rect 412270 117399 412326 117408
rect 412180 57928 412232 57934
rect 412180 57870 412232 57876
rect 412178 56536 412234 56545
rect 412178 56471 412234 56480
rect 412192 40730 412220 56471
rect 412284 46918 412312 117399
rect 412362 97880 412418 97889
rect 412362 97815 412418 97824
rect 412272 46912 412324 46918
rect 412272 46854 412324 46860
rect 412270 44840 412326 44849
rect 412270 44775 412326 44784
rect 412180 40724 412232 40730
rect 412180 40666 412232 40672
rect 412088 33040 412140 33046
rect 412088 32982 412140 32988
rect 412284 31754 412312 44775
rect 412272 31748 412324 31754
rect 412272 31690 412324 31696
rect 412376 31618 412404 97815
rect 412468 93854 412496 128318
rect 412468 93826 412588 93854
rect 412560 80209 412588 93826
rect 412546 80200 412602 80209
rect 412546 80135 412602 80144
rect 413296 64530 413324 129950
rect 413468 129940 413520 129946
rect 413468 129882 413520 129888
rect 413376 129804 413428 129810
rect 413376 129746 413428 129752
rect 413388 93974 413416 129746
rect 413376 93968 413428 93974
rect 413376 93910 413428 93916
rect 413376 89820 413428 89826
rect 413376 89762 413428 89768
rect 413284 64524 413336 64530
rect 413284 64466 413336 64472
rect 413284 52556 413336 52562
rect 413284 52498 413336 52504
rect 412454 50688 412510 50697
rect 412454 50623 412510 50632
rect 412364 31612 412416 31618
rect 412364 31554 412416 31560
rect 411904 30184 411956 30190
rect 411904 30126 411956 30132
rect 412468 30122 412496 50623
rect 412546 46744 412602 46753
rect 412546 46679 412602 46688
rect 412560 31686 412588 46679
rect 412548 31680 412600 31686
rect 412548 31622 412600 31628
rect 412456 30116 412508 30122
rect 412456 30058 412508 30064
rect 410616 29300 410668 29306
rect 410616 29242 410668 29248
rect 410524 29232 410576 29238
rect 410524 29174 410576 29180
rect 405738 28928 405794 28937
rect 405738 28863 405794 28872
rect 389180 28766 389232 28772
rect 397458 28792 397514 28801
rect 356612 28756 356664 28762
rect 397458 28727 397514 28736
rect 356612 28698 356664 28704
rect 348516 28688 348568 28694
rect 348516 28630 348568 28636
rect 413296 28626 413324 52498
rect 413388 28966 413416 89762
rect 413480 76770 413508 129882
rect 413836 127016 413888 127022
rect 413836 126958 413888 126964
rect 413744 125656 413796 125662
rect 413744 125598 413796 125604
rect 413652 124228 413704 124234
rect 413652 124170 413704 124176
rect 413560 122868 413612 122874
rect 413560 122810 413612 122816
rect 413468 76764 413520 76770
rect 413468 76706 413520 76712
rect 413572 74254 413600 122810
rect 413664 78266 413692 124170
rect 413756 84182 413784 125598
rect 413848 86494 413876 126958
rect 413836 86488 413888 86494
rect 413836 86430 413888 86436
rect 413744 84176 413796 84182
rect 413744 84118 413796 84124
rect 413652 78260 413704 78266
rect 413652 78202 413704 78208
rect 413560 74248 413612 74254
rect 413560 74190 413612 74196
rect 413468 54052 413520 54058
rect 413468 53994 413520 54000
rect 413480 29306 413508 53994
rect 414676 38894 414704 131310
rect 414756 131300 414808 131306
rect 414756 131242 414808 131248
rect 414768 41070 414796 131242
rect 414848 131232 414900 131238
rect 414848 131174 414900 131180
rect 414860 42702 414888 131174
rect 414952 74526 414980 151778
rect 415032 147688 415084 147694
rect 415032 147630 415084 147636
rect 414940 74520 414992 74526
rect 414940 74462 414992 74468
rect 415044 71738 415072 147630
rect 415216 129872 415268 129878
rect 415216 129814 415268 129820
rect 415124 100768 415176 100774
rect 415124 100710 415176 100716
rect 415032 71732 415084 71738
rect 415032 71674 415084 71680
rect 414848 42696 414900 42702
rect 414848 42638 414900 42644
rect 414756 41064 414808 41070
rect 414756 41006 414808 41012
rect 414664 38888 414716 38894
rect 414664 38830 414716 38836
rect 415136 34474 415164 100710
rect 415228 95878 415256 129814
rect 416056 109002 416084 195978
rect 416136 184952 416188 184958
rect 416136 184894 416188 184900
rect 416044 108996 416096 109002
rect 416044 108938 416096 108944
rect 416044 103556 416096 103562
rect 416044 103498 416096 103504
rect 415216 95872 415268 95878
rect 415216 95814 415268 95820
rect 416056 35902 416084 103498
rect 416148 102134 416176 184894
rect 417424 165640 417476 165646
rect 417424 165582 417476 165588
rect 416228 124296 416280 124302
rect 416228 124238 416280 124244
rect 416136 102128 416188 102134
rect 416136 102070 416188 102076
rect 416240 53786 416268 124238
rect 416320 118720 416372 118726
rect 416320 118662 416372 118668
rect 416228 53780 416280 53786
rect 416228 53722 416280 53728
rect 416332 48278 416360 118662
rect 416412 113212 416464 113218
rect 416412 113154 416464 113160
rect 416320 48272 416372 48278
rect 416320 48214 416372 48220
rect 416424 44130 416452 113154
rect 416504 107704 416556 107710
rect 416504 107646 416556 107652
rect 416412 44124 416464 44130
rect 416412 44066 416464 44072
rect 416516 38622 416544 107646
rect 417436 85542 417464 165582
rect 417608 161492 417660 161498
rect 417608 161434 417660 161440
rect 417516 158772 417568 158778
rect 417516 158714 417568 158720
rect 417424 85536 417476 85542
rect 417424 85478 417476 85484
rect 417528 80034 417556 158714
rect 417620 82822 417648 161434
rect 417700 154624 417752 154630
rect 417700 154566 417752 154572
rect 417608 82816 417660 82822
rect 417608 82758 417660 82764
rect 417516 80028 417568 80034
rect 417516 79970 417568 79976
rect 417712 77246 417740 154566
rect 417792 150476 417844 150482
rect 417792 150418 417844 150424
rect 417700 77240 417752 77246
rect 417700 77182 417752 77188
rect 417804 73098 417832 150418
rect 417884 144968 417936 144974
rect 417884 144910 417936 144916
rect 417792 73092 417844 73098
rect 417792 73034 417844 73040
rect 417896 68950 417924 144910
rect 417976 109064 418028 109070
rect 417976 109006 418028 109012
rect 417884 68944 417936 68950
rect 417884 68886 417936 68892
rect 417424 59424 417476 59430
rect 417424 59366 417476 59372
rect 416504 38616 416556 38622
rect 416504 38558 416556 38564
rect 416044 35896 416096 35902
rect 416044 35838 416096 35844
rect 415124 34468 415176 34474
rect 415124 34410 415176 34416
rect 413468 29300 413520 29306
rect 413468 29242 413520 29248
rect 413376 28960 413428 28966
rect 413376 28902 413428 28908
rect 417436 28762 417464 59366
rect 417516 48340 417568 48346
rect 417516 48282 417568 48288
rect 417528 29374 417556 48282
rect 417988 41410 418016 109006
rect 417976 41404 418028 41410
rect 417976 41346 418028 41352
rect 417516 29368 417568 29374
rect 417516 29310 417568 29316
rect 417424 28756 417476 28762
rect 417424 28698 417476 28704
rect 340420 28620 340472 28626
rect 340420 28562 340472 28568
rect 413284 28620 413336 28626
rect 413284 28562 413336 28568
rect 332140 28552 332192 28558
rect 332140 28494 332192 28500
rect 324412 28484 324464 28490
rect 324412 28426 324464 28432
rect 316132 28416 316184 28422
rect 316132 28358 316184 28364
rect 307760 28348 307812 28354
rect 307760 28290 307812 28296
rect 283380 28280 283432 28286
rect 283380 28222 283432 28228
rect 275100 28212 275152 28218
rect 275100 28154 275152 28160
rect 267004 28144 267056 28150
rect 267004 28086 267056 28092
rect 234620 28076 234672 28082
rect 234620 28018 234672 28024
rect 418816 20670 418844 209782
rect 421564 197396 421616 197402
rect 421564 197338 421616 197344
rect 418988 169788 419040 169794
rect 418988 169730 419040 169736
rect 418896 130076 418948 130082
rect 418896 130018 418948 130024
rect 418908 35834 418936 130018
rect 419000 89690 419028 169730
rect 420276 168428 420328 168434
rect 420276 168370 420328 168376
rect 420184 164280 420236 164286
rect 420184 164222 420236 164228
rect 419080 155984 419132 155990
rect 419080 155926 419132 155932
rect 418988 89684 419040 89690
rect 418988 89626 419040 89632
rect 419092 78674 419120 155926
rect 419356 131504 419408 131510
rect 419356 131446 419408 131452
rect 419264 128444 419316 128450
rect 419264 128386 419316 128392
rect 419172 114572 419224 114578
rect 419172 114514 419224 114520
rect 419080 78668 419132 78674
rect 419080 78610 419132 78616
rect 418988 69080 419040 69086
rect 418988 69022 419040 69028
rect 418896 35828 418948 35834
rect 418896 35770 418948 35776
rect 419000 28898 419028 69022
rect 419184 45558 419212 114514
rect 419276 88330 419304 128386
rect 419368 92478 419396 131446
rect 419356 92472 419408 92478
rect 419356 92414 419408 92420
rect 419264 88324 419316 88330
rect 419264 88266 419316 88272
rect 420196 84182 420224 164222
rect 420288 88330 420316 168370
rect 420368 160132 420420 160138
rect 420368 160074 420420 160080
rect 420276 88324 420328 88330
rect 420276 88266 420328 88272
rect 420184 84176 420236 84182
rect 420184 84118 420236 84124
rect 420380 81394 420408 160074
rect 420460 132524 420512 132530
rect 420460 132466 420512 132472
rect 420368 81388 420420 81394
rect 420368 81330 420420 81336
rect 420472 59362 420500 132466
rect 420552 128512 420604 128518
rect 420552 128454 420604 128460
rect 420460 59356 420512 59362
rect 420460 59298 420512 59304
rect 420564 56574 420592 128454
rect 421576 110430 421604 197338
rect 436744 191888 436796 191894
rect 436744 191830 436796 191836
rect 421656 189100 421708 189106
rect 421656 189042 421708 189048
rect 421564 110424 421616 110430
rect 421564 110366 421616 110372
rect 421668 104854 421696 189042
rect 435364 187740 435416 187746
rect 435364 187682 435416 187688
rect 432604 183592 432656 183598
rect 432604 183534 432656 183540
rect 431224 182232 431276 182238
rect 431224 182174 431276 182180
rect 429844 179444 429896 179450
rect 429844 179386 429896 179392
rect 428464 178084 428516 178090
rect 428464 178026 428516 178032
rect 425704 175296 425756 175302
rect 425704 175238 425756 175244
rect 424324 173936 424376 173942
rect 424324 173878 424376 173884
rect 421748 172576 421800 172582
rect 421748 172518 421800 172524
rect 421656 104848 421708 104854
rect 421656 104790 421708 104796
rect 421760 91050 421788 172518
rect 421840 146328 421892 146334
rect 421840 146270 421892 146276
rect 421748 91044 421800 91050
rect 421748 90986 421800 90992
rect 421852 70378 421880 146270
rect 421932 140820 421984 140826
rect 421932 140762 421984 140768
rect 421840 70372 421892 70378
rect 421840 70314 421892 70320
rect 421944 66230 421972 140762
rect 422024 136672 422076 136678
rect 422024 136614 422076 136620
rect 421932 66224 421984 66230
rect 421932 66166 421984 66172
rect 422036 62082 422064 136614
rect 423772 121576 423824 121582
rect 423772 121518 423824 121524
rect 423784 120766 423812 121518
rect 423772 120760 423824 120766
rect 423772 120702 423824 120708
rect 424336 92478 424364 173878
rect 425716 93838 425744 175238
rect 425796 128512 425848 128518
rect 425796 128454 425848 128460
rect 425808 121582 425836 128454
rect 425796 121576 425848 121582
rect 425796 121518 425848 121524
rect 428476 95198 428504 178026
rect 428556 122936 428608 122942
rect 428556 122878 428608 122884
rect 428464 95192 428516 95198
rect 428464 95134 428516 95140
rect 425704 93832 425756 93838
rect 425704 93774 425756 93780
rect 424324 92472 424376 92478
rect 424324 92414 424376 92420
rect 422024 62076 422076 62082
rect 422024 62018 422076 62024
rect 420552 56568 420604 56574
rect 420552 56510 420604 56516
rect 428568 52426 428596 122878
rect 429856 96626 429884 179386
rect 429936 142180 429988 142186
rect 429936 142122 429988 142128
rect 429844 96620 429896 96626
rect 429844 96562 429896 96568
rect 429948 67590 429976 142122
rect 431236 97986 431264 182174
rect 431316 138032 431368 138038
rect 431316 137974 431368 137980
rect 431224 97980 431276 97986
rect 431224 97922 431276 97928
rect 429936 67584 429988 67590
rect 429936 67526 429988 67532
rect 431328 64870 431356 137974
rect 432616 100706 432644 183534
rect 432696 133952 432748 133958
rect 432696 133894 432748 133900
rect 432604 100700 432656 100706
rect 432604 100642 432656 100648
rect 431316 64864 431368 64870
rect 431316 64806 431368 64812
rect 432708 60722 432736 133894
rect 434628 130416 434680 130422
rect 434628 130358 434680 130364
rect 434640 128518 434668 130358
rect 434628 128512 434680 128518
rect 434628 128454 434680 128460
rect 435376 103086 435404 187682
rect 435456 127084 435508 127090
rect 435456 127026 435508 127032
rect 435364 103080 435416 103086
rect 435364 103022 435416 103028
rect 432696 60716 432748 60722
rect 432696 60658 432748 60664
rect 435468 54738 435496 127026
rect 436756 106185 436784 191830
rect 463712 151814 463740 231814
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218074 580212 218991
rect 543004 218068 543056 218074
rect 543004 218010 543056 218016
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 540244 202904 540296 202910
rect 540244 202846 540296 202852
rect 463712 151786 464568 151814
rect 444656 131436 444708 131442
rect 444656 131378 444708 131384
rect 444668 129962 444696 131378
rect 454592 130416 454644 130422
rect 454592 130358 454644 130364
rect 454604 129962 454632 130358
rect 464540 129962 464568 151786
rect 534632 131504 534684 131510
rect 534632 131446 534684 131452
rect 484584 131368 484636 131374
rect 484584 131310 484636 131316
rect 474740 130076 474792 130082
rect 474740 130018 474792 130024
rect 474752 129962 474780 130018
rect 484596 129962 484624 131310
rect 494612 131300 494664 131306
rect 494612 131242 494664 131248
rect 494624 129962 494652 131242
rect 504640 131232 504692 131238
rect 504640 131174 504692 131180
rect 504652 129962 504680 131174
rect 514760 130008 514812 130014
rect 444668 129934 445004 129962
rect 454604 129934 454940 129962
rect 464540 129934 464968 129962
rect 474752 129934 474996 129962
rect 484596 129934 484932 129962
rect 494624 129934 494960 129962
rect 504652 129934 504988 129962
rect 534644 129962 534672 131446
rect 514812 129956 514924 129962
rect 514760 129950 514924 129956
rect 514772 129934 514924 129950
rect 524616 129946 524952 129962
rect 524604 129940 524952 129946
rect 524656 129934 524952 129940
rect 534644 129934 534980 129962
rect 524604 129882 524656 129888
rect 539324 129872 539376 129878
rect 539324 129814 539376 129820
rect 437478 128752 437534 128761
rect 437478 128687 437534 128696
rect 437492 128450 437520 128687
rect 437480 128444 437532 128450
rect 437480 128386 437532 128392
rect 437478 127392 437534 127401
rect 437478 127327 437534 127336
rect 437492 127022 437520 127327
rect 437480 127016 437532 127022
rect 437480 126958 437532 126964
rect 539336 126041 539364 129814
rect 539322 126032 539378 126041
rect 539322 125967 539378 125976
rect 437478 125896 437534 125905
rect 437478 125831 437534 125840
rect 437492 125662 437520 125831
rect 437480 125656 437532 125662
rect 437480 125598 437532 125604
rect 437478 124264 437534 124273
rect 437478 124199 437480 124208
rect 437532 124199 437534 124208
rect 437480 124170 437532 124176
rect 437478 123040 437534 123049
rect 437478 122975 437534 122984
rect 437492 122874 437520 122975
rect 437480 122868 437532 122874
rect 437480 122810 437532 122816
rect 438490 120864 438546 120873
rect 438490 120799 438546 120808
rect 436836 120148 436888 120154
rect 436836 120090 436888 120096
rect 436742 106176 436798 106185
rect 436742 106111 436798 106120
rect 436744 66292 436796 66298
rect 436744 66234 436796 66240
rect 435456 54732 435508 54738
rect 435456 54674 435508 54680
rect 428556 52420 428608 52426
rect 428556 52362 428608 52368
rect 419172 45552 419224 45558
rect 419172 45494 419224 45500
rect 418988 28892 419040 28898
rect 418988 28834 419040 28840
rect 436756 28694 436784 66234
rect 436848 49609 436876 120090
rect 438398 119232 438454 119241
rect 438398 119167 438454 119176
rect 438306 117736 438362 117745
rect 438306 117671 438362 117680
rect 438214 116104 438270 116113
rect 438214 116039 438270 116048
rect 438122 114608 438178 114617
rect 438122 114543 438178 114552
rect 437480 114504 437532 114510
rect 437480 114446 437532 114452
rect 437492 114073 437520 114446
rect 437478 114064 437534 114073
rect 437478 113999 437534 114008
rect 437480 113144 437532 113150
rect 437480 113086 437532 113092
rect 437492 112577 437520 113086
rect 437478 112568 437534 112577
rect 437478 112503 437534 112512
rect 437480 110424 437532 110430
rect 437480 110366 437532 110372
rect 437492 110265 437520 110366
rect 437478 110256 437534 110265
rect 437478 110191 437534 110200
rect 437478 109032 437534 109041
rect 437478 108967 437480 108976
rect 437532 108967 437534 108976
rect 437480 108938 437532 108944
rect 437480 107636 437532 107642
rect 437480 107578 437532 107584
rect 437492 107409 437520 107578
rect 437478 107400 437534 107409
rect 437478 107335 437534 107344
rect 437480 104848 437532 104854
rect 437480 104790 437532 104796
rect 437492 104553 437520 104790
rect 437478 104544 437534 104553
rect 437478 104479 437534 104488
rect 437664 103080 437716 103086
rect 437662 103048 437664 103057
rect 437716 103048 437718 103057
rect 437662 102983 437718 102992
rect 437480 102128 437532 102134
rect 437480 102070 437532 102076
rect 437492 101561 437520 102070
rect 437478 101552 437534 101561
rect 437478 101487 437534 101496
rect 437480 100700 437532 100706
rect 437480 100642 437532 100648
rect 437492 100065 437520 100642
rect 437478 100056 437534 100065
rect 437478 99991 437534 100000
rect 437480 97980 437532 97986
rect 437480 97922 437532 97928
rect 437492 97753 437520 97922
rect 437478 97744 437534 97753
rect 437478 97679 437534 97688
rect 437480 96620 437532 96626
rect 437480 96562 437532 96568
rect 437492 96529 437520 96562
rect 437478 96520 437534 96529
rect 437478 96455 437534 96464
rect 437480 95192 437532 95198
rect 437478 95160 437480 95169
rect 437532 95160 437534 95169
rect 437478 95095 437534 95104
rect 437480 93832 437532 93838
rect 437480 93774 437532 93780
rect 437492 93537 437520 93774
rect 437478 93528 437534 93537
rect 437478 93463 437534 93472
rect 437480 92472 437532 92478
rect 437480 92414 437532 92420
rect 437492 92041 437520 92414
rect 437478 92032 437534 92041
rect 437478 91967 437534 91976
rect 437480 91044 437532 91050
rect 437480 90986 437532 90992
rect 437492 90545 437520 90986
rect 437478 90536 437534 90545
rect 437478 90471 437534 90480
rect 437480 89684 437532 89690
rect 437480 89626 437532 89632
rect 437492 89049 437520 89626
rect 437478 89040 437534 89049
rect 437478 88975 437534 88984
rect 437480 88324 437532 88330
rect 437480 88266 437532 88272
rect 437492 87553 437520 88266
rect 437478 87544 437534 87553
rect 437478 87479 437534 87488
rect 437480 85536 437532 85542
rect 437478 85504 437480 85513
rect 437532 85504 437534 85513
rect 437478 85439 437534 85448
rect 437480 84176 437532 84182
rect 437478 84144 437480 84153
rect 437532 84144 437534 84153
rect 437478 84079 437534 84088
rect 437480 82816 437532 82822
rect 437480 82758 437532 82764
rect 437492 82521 437520 82758
rect 437478 82512 437534 82521
rect 437478 82447 437534 82456
rect 437480 81388 437532 81394
rect 437480 81330 437532 81336
rect 437492 81025 437520 81330
rect 437478 81016 437534 81025
rect 437478 80951 437534 80960
rect 437480 80028 437532 80034
rect 437480 79970 437532 79976
rect 437492 79665 437520 79970
rect 437478 79656 437534 79665
rect 437478 79591 437534 79600
rect 437480 78668 437532 78674
rect 437480 78610 437532 78616
rect 437492 78169 437520 78610
rect 437478 78160 437534 78169
rect 437478 78095 437534 78104
rect 437480 77240 437532 77246
rect 437480 77182 437532 77188
rect 437492 76673 437520 77182
rect 437478 76664 437534 76673
rect 437478 76599 437534 76608
rect 437480 74520 437532 74526
rect 437480 74462 437532 74468
rect 437492 74361 437520 74462
rect 437478 74352 437534 74361
rect 437478 74287 437534 74296
rect 437478 73128 437534 73137
rect 437478 73063 437480 73072
rect 437532 73063 437534 73072
rect 437480 73034 437532 73040
rect 437480 71732 437532 71738
rect 437480 71674 437532 71680
rect 437492 71505 437520 71674
rect 437478 71496 437534 71505
rect 437478 71431 437534 71440
rect 437480 70372 437532 70378
rect 437480 70314 437532 70320
rect 437492 70281 437520 70314
rect 437478 70272 437534 70281
rect 437478 70207 437534 70216
rect 437480 68944 437532 68950
rect 437480 68886 437532 68892
rect 437492 68649 437520 68886
rect 437478 68640 437534 68649
rect 437478 68575 437534 68584
rect 437480 67584 437532 67590
rect 437480 67526 437532 67532
rect 437492 67153 437520 67526
rect 437478 67144 437534 67153
rect 437478 67079 437534 67088
rect 437480 66224 437532 66230
rect 437480 66166 437532 66172
rect 437492 65657 437520 66166
rect 437478 65648 437534 65657
rect 437478 65583 437534 65592
rect 437480 64864 437532 64870
rect 437480 64806 437532 64812
rect 437492 64161 437520 64806
rect 437478 64152 437534 64161
rect 437478 64087 437534 64096
rect 437478 62112 437534 62121
rect 437478 62047 437480 62056
rect 437532 62047 437534 62056
rect 437480 62018 437532 62024
rect 437480 60716 437532 60722
rect 437480 60658 437532 60664
rect 437492 60625 437520 60658
rect 437478 60616 437534 60625
rect 437478 60551 437534 60560
rect 437480 59356 437532 59362
rect 437480 59298 437532 59304
rect 437492 59265 437520 59298
rect 437478 59256 437534 59265
rect 437478 59191 437534 59200
rect 437480 57928 437532 57934
rect 437480 57870 437532 57876
rect 437492 57633 437520 57870
rect 437478 57624 437534 57633
rect 437478 57559 437534 57568
rect 437480 56568 437532 56574
rect 437480 56510 437532 56516
rect 437492 56137 437520 56510
rect 437478 56128 437534 56137
rect 437478 56063 437534 56072
rect 437756 54732 437808 54738
rect 437756 54674 437808 54680
rect 437768 54641 437796 54674
rect 437754 54632 437810 54641
rect 437754 54567 437810 54576
rect 437480 53780 437532 53786
rect 437480 53722 437532 53728
rect 437492 53145 437520 53722
rect 437478 53136 437534 53145
rect 437478 53071 437534 53080
rect 437480 52420 437532 52426
rect 437480 52362 437532 52368
rect 437492 51649 437520 52362
rect 437478 51640 437534 51649
rect 437478 51575 437534 51584
rect 436834 49600 436890 49609
rect 436834 49535 436890 49544
rect 437480 48272 437532 48278
rect 437478 48240 437480 48249
rect 437532 48240 437534 48249
rect 437478 48175 437534 48184
rect 437480 46912 437532 46918
rect 437480 46854 437532 46860
rect 437492 46617 437520 46854
rect 437478 46608 437534 46617
rect 437478 46543 437534 46552
rect 437480 45552 437532 45558
rect 437480 45494 437532 45500
rect 437492 45257 437520 45494
rect 437478 45248 437534 45257
rect 437478 45183 437534 45192
rect 437480 44124 437532 44130
rect 437480 44066 437532 44072
rect 437492 43625 437520 44066
rect 437478 43616 437534 43625
rect 437478 43551 437534 43560
rect 437480 42764 437532 42770
rect 437480 42706 437532 42712
rect 437492 42265 437520 42706
rect 437478 42256 437534 42265
rect 437478 42191 437534 42200
rect 437480 41404 437532 41410
rect 437480 41346 437532 41352
rect 437492 40633 437520 41346
rect 437478 40624 437534 40633
rect 437478 40559 437534 40568
rect 437480 38616 437532 38622
rect 437480 38558 437532 38564
rect 437492 38457 437520 38558
rect 437478 38448 437534 38457
rect 437478 38383 437534 38392
rect 437480 37256 437532 37262
rect 437478 37224 437480 37233
rect 437532 37224 437534 37233
rect 437478 37159 437534 37168
rect 437480 35896 437532 35902
rect 437478 35864 437480 35873
rect 437532 35864 437534 35873
rect 437478 35799 437534 35808
rect 437480 34468 437532 34474
rect 437480 34410 437532 34416
rect 437492 34105 437520 34410
rect 437478 34096 437534 34105
rect 437478 34031 437534 34040
rect 438136 33114 438164 114543
rect 438228 37194 438256 116039
rect 438320 63510 438348 117671
rect 438412 69018 438440 119167
rect 438504 73166 438532 120799
rect 540256 100706 540284 202846
rect 542452 129804 542504 129810
rect 542452 129746 542504 129752
rect 542360 128376 542412 128382
rect 542360 128318 542412 128324
rect 542372 107273 542400 128318
rect 542464 116385 542492 129746
rect 542450 116376 542506 116385
rect 542450 116311 542506 116320
rect 542358 107264 542414 107273
rect 542358 107199 542414 107208
rect 540244 100700 540296 100706
rect 540244 100642 540296 100648
rect 542358 98152 542414 98161
rect 542358 98087 542414 98096
rect 439504 81456 439556 81462
rect 439504 81398 439556 81404
rect 438492 73160 438544 73166
rect 438492 73102 438544 73108
rect 438400 69012 438452 69018
rect 438400 68954 438452 68960
rect 438308 63504 438360 63510
rect 438308 63446 438360 63452
rect 438216 37188 438268 37194
rect 438216 37130 438268 37136
rect 438124 33108 438176 33114
rect 438124 33050 438176 33056
rect 437480 33040 437532 33046
rect 437480 32982 437532 32988
rect 437492 32745 437520 32982
rect 437478 32736 437534 32745
rect 437478 32671 437534 32680
rect 437480 31612 437532 31618
rect 437480 31554 437532 31560
rect 437492 31249 437520 31554
rect 437478 31240 437534 31249
rect 437478 31175 437534 31184
rect 439516 28830 439544 81398
rect 439596 57996 439648 58002
rect 439596 57938 439648 57944
rect 439504 28824 439556 28830
rect 439504 28766 439556 28772
rect 436744 28688 436796 28694
rect 436744 28630 436796 28636
rect 439608 28558 439636 57938
rect 542372 30190 542400 98087
rect 542450 89040 542506 89049
rect 542450 88975 542506 88984
rect 542360 30184 542412 30190
rect 444176 30110 444328 30138
rect 452456 30110 452608 30138
rect 444300 29170 444328 30110
rect 452580 29238 452608 30110
rect 460492 30110 460828 30138
rect 468772 30110 469108 30138
rect 477480 30110 477540 30138
rect 485760 30110 485820 30138
rect 494132 30110 494192 30138
rect 452568 29232 452620 29238
rect 452568 29174 452620 29180
rect 444288 29164 444340 29170
rect 444288 29106 444340 29112
rect 439596 28552 439648 28558
rect 439596 28494 439648 28500
rect 460492 27606 460520 30110
rect 468772 29374 468800 30110
rect 468760 29368 468812 29374
rect 468760 29310 468812 29316
rect 477512 28626 477540 30110
rect 485792 29306 485820 30110
rect 485780 29300 485832 29306
rect 485780 29242 485832 29248
rect 477500 28620 477552 28626
rect 477500 28562 477552 28568
rect 494164 28558 494192 30110
rect 502352 30110 502504 30138
rect 510632 30110 510784 30138
rect 519004 30110 519156 30138
rect 527192 30110 527436 30138
rect 535472 30110 535808 30138
rect 542360 30126 542412 30132
rect 542464 30122 542492 88975
rect 542542 80064 542598 80073
rect 542542 79999 542598 80008
rect 542556 31686 542584 79999
rect 542634 70952 542690 70961
rect 542634 70887 542690 70896
rect 542648 31754 542676 70887
rect 542726 61840 542782 61849
rect 542726 61775 542782 61784
rect 542636 31748 542688 31754
rect 542636 31690 542688 31696
rect 542544 31680 542596 31686
rect 542544 31622 542596 31628
rect 542740 30258 542768 61775
rect 543016 43625 543044 218010
rect 544384 205692 544436 205698
rect 544384 205634 544436 205640
rect 543188 191888 543240 191894
rect 543188 191830 543240 191836
rect 543096 178084 543148 178090
rect 543096 178026 543148 178032
rect 543002 43616 543058 43625
rect 543002 43551 543058 43560
rect 543108 34649 543136 178026
rect 543200 52737 543228 191830
rect 544396 60722 544424 205634
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580184 191894 580212 192471
rect 580172 191888 580224 191894
rect 580172 191830 580224 191836
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580276 112849 580304 248406
rect 580368 152697 580396 249766
rect 580354 152688 580410 152697
rect 580354 152623 580410 152632
rect 580354 126032 580410 126041
rect 580354 125967 580410 125976
rect 580262 112840 580318 112849
rect 580262 112775 580318 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580262 86184 580318 86193
rect 580262 86119 580318 86128
rect 544384 60716 544436 60722
rect 544384 60658 544436 60664
rect 579804 60716 579856 60722
rect 579804 60658 579856 60664
rect 579816 59673 579844 60658
rect 579802 59664 579858 59673
rect 579802 59599 579858 59608
rect 543186 52728 543242 52737
rect 543186 52663 543242 52672
rect 543094 34640 543150 34649
rect 543094 34575 543150 34584
rect 580170 33144 580226 33153
rect 580170 33079 580226 33088
rect 580184 30326 580212 33079
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 542728 30252 542780 30258
rect 542728 30194 542780 30200
rect 542452 30116 542504 30122
rect 502352 28762 502380 30110
rect 502340 28756 502392 28762
rect 502340 28698 502392 28704
rect 510632 28694 510660 30110
rect 519004 28898 519032 30110
rect 518992 28892 519044 28898
rect 518992 28834 519044 28840
rect 527192 28830 527220 30110
rect 535472 28966 535500 30110
rect 542452 30058 542504 30064
rect 580276 29170 580304 86119
rect 580368 29238 580396 125967
rect 580446 72992 580502 73001
rect 580446 72927 580502 72936
rect 580356 29232 580408 29238
rect 580356 29174 580408 29180
rect 580264 29164 580316 29170
rect 580264 29106 580316 29112
rect 580460 29102 580488 72927
rect 580538 46336 580594 46345
rect 580538 46271 580594 46280
rect 580448 29096 580500 29102
rect 580448 29038 580500 29044
rect 580552 29034 580580 46271
rect 580540 29028 580592 29034
rect 580540 28970 580592 28976
rect 535460 28960 535512 28966
rect 535460 28902 535512 28908
rect 527180 28824 527232 28830
rect 527180 28766 527232 28772
rect 510620 28688 510672 28694
rect 510620 28630 510672 28636
rect 494152 28552 494204 28558
rect 494152 28494 494204 28500
rect 460480 27600 460532 27606
rect 460480 27542 460532 27548
rect 418804 20664 418856 20670
rect 418804 20606 418856 20612
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 218060 6860 218112 6866
rect 218060 6802 218112 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 201500 4140 201552 4146
rect 201500 4082 201552 4088
rect 193220 4072 193272 4078
rect 193220 4014 193272 4020
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 572 3664 624 3670
rect 572 3606 624 3612
rect 1308 3664 1360 3670
rect 1308 3606 1360 3612
rect 584 480 612 3606
rect 1688 480 1716 3674
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 48226 334192 48282 334248
rect 48134 332968 48190 333024
rect 47950 331064 48006 331120
rect 47858 328480 47914 328536
rect 47766 327528 47822 327584
rect 47674 305632 47730 305688
rect 48042 325760 48098 325816
rect 208306 334056 208362 334112
rect 49606 330066 49662 330122
rect 49514 307218 49570 307274
rect 208214 329976 208270 330032
rect 208122 328480 208178 328536
rect 208030 327392 208086 327448
rect 207018 325760 207074 325816
rect 55862 299512 55918 299568
rect 103242 298152 103298 298208
rect 65706 298016 65762 298072
rect 67546 298016 67602 298072
rect 67822 298016 67878 298072
rect 69938 298016 69994 298072
rect 70214 298016 70270 298072
rect 71502 298016 71558 298072
rect 73066 298016 73122 298072
rect 74446 298016 74502 298072
rect 75826 298016 75882 298072
rect 76838 298016 76894 298072
rect 77114 298016 77170 298072
rect 78586 298016 78642 298072
rect 79874 298016 79930 298072
rect 81254 298016 81310 298072
rect 81806 298016 81862 298072
rect 82634 298016 82690 298072
rect 84014 298016 84070 298072
rect 85302 298016 85358 298072
rect 86774 298016 86830 298072
rect 88154 298016 88210 298072
rect 89626 298016 89682 298072
rect 90914 298016 90970 298072
rect 92386 298016 92442 298072
rect 93306 298016 93362 298072
rect 93674 298016 93730 298072
rect 95054 298016 95110 298072
rect 96526 298016 96582 298072
rect 96710 298016 96766 298072
rect 97814 298016 97870 298072
rect 99286 298016 99342 298072
rect 100574 298016 100630 298072
rect 101862 298016 101918 298072
rect 78494 297880 78550 297936
rect 79782 297880 79838 297936
rect 81346 297880 81402 297936
rect 84106 297880 84162 297936
rect 85394 297880 85450 297936
rect 86682 297880 86738 297936
rect 85486 297064 85542 297120
rect 86866 297744 86922 297800
rect 88246 297880 88302 297936
rect 89534 297880 89590 297936
rect 91006 297880 91062 297936
rect 92294 297880 92350 297936
rect 93582 297880 93638 297936
rect 95146 297880 95202 297936
rect 96434 297880 96490 297936
rect 97722 297880 97778 297936
rect 99194 297880 99250 297936
rect 100666 297880 100722 297936
rect 102046 297880 102102 297936
rect 101954 297744 102010 297800
rect 103334 298016 103390 298072
rect 104806 298016 104862 298072
rect 106186 298016 106242 298072
rect 106738 298016 106794 298072
rect 107474 298016 107530 298072
rect 108946 298016 109002 298072
rect 110326 298016 110382 298072
rect 111706 298016 111762 298072
rect 112994 298016 113050 298072
rect 114466 298016 114522 298072
rect 115846 298016 115902 298072
rect 117226 298016 117282 298072
rect 104714 297880 104770 297936
rect 106094 297880 106150 297936
rect 108854 297880 108910 297936
rect 113086 297880 113142 297936
rect 187606 249464 187662 249520
rect 187330 246064 187386 246120
rect 187514 248376 187570 248432
rect 187606 247288 187662 247344
rect 187606 244976 187662 245032
rect 186318 243888 186374 243944
rect 186318 242664 186374 242720
rect 186410 241576 186466 241632
rect 186318 240488 186374 240544
rect 186318 239400 186374 239456
rect 186318 238176 186374 238232
rect 186318 237088 186374 237144
rect 186410 236000 186466 236056
rect 186318 234776 186374 234832
rect 186318 233688 186374 233744
rect 186318 232600 186374 232656
rect 186318 231376 186374 231432
rect 186318 229200 186374 229256
rect 186318 228112 186374 228168
rect 186686 225664 186742 225720
rect 186318 222264 186374 222320
rect 131118 129684 131120 129704
rect 131120 129684 131172 129704
rect 131172 129684 131174 129704
rect 131118 129648 131174 129684
rect 131210 128560 131266 128616
rect 131210 127336 131266 127392
rect 131210 126828 131212 126848
rect 131212 126828 131264 126848
rect 131264 126828 131266 126848
rect 131210 126792 131266 126828
rect 131118 126112 131174 126168
rect 131118 125568 131174 125624
rect 131578 125024 131634 125080
rect 131210 124480 131266 124536
rect 131118 123256 131174 123312
rect 131854 129104 131910 129160
rect 131762 127880 131818 127936
rect 131762 123800 131818 123856
rect 131210 122732 131266 122768
rect 131210 122712 131212 122732
rect 131212 122712 131264 122732
rect 131264 122712 131266 122732
rect 131486 122032 131542 122088
rect 131118 121488 131174 121544
rect 131210 120944 131266 121000
rect 131118 120264 131174 120320
rect 131118 119176 131174 119232
rect 131210 118532 131212 118552
rect 131212 118532 131264 118552
rect 131264 118532 131266 118552
rect 131210 118496 131266 118532
rect 131302 117952 131358 118008
rect 131118 117408 131174 117464
rect 131210 116864 131266 116920
rect 131118 116184 131174 116240
rect 131210 115096 131266 115152
rect 131210 114436 131266 114472
rect 131210 114416 131212 114436
rect 131212 114416 131264 114436
rect 131264 114416 131266 114436
rect 131118 113872 131174 113928
rect 131302 113328 131358 113384
rect 131210 112784 131266 112840
rect 131118 112104 131174 112160
rect 131210 111560 131266 111616
rect 131118 111016 131174 111072
rect 131210 110372 131212 110392
rect 131212 110372 131264 110392
rect 131264 110372 131266 110392
rect 131210 110336 131266 110372
rect 131210 109792 131266 109848
rect 131118 109248 131174 109304
rect 131210 108568 131266 108624
rect 131118 108024 131174 108080
rect 131210 107500 131266 107536
rect 131210 107480 131212 107500
rect 131212 107480 131264 107500
rect 131264 107480 131266 107500
rect 131118 106936 131174 106992
rect 131302 106256 131358 106312
rect 131210 105712 131266 105768
rect 131118 105168 131174 105224
rect 131210 104488 131266 104544
rect 131118 103944 131174 104000
rect 131210 103420 131266 103456
rect 131210 103400 131212 103420
rect 131212 103400 131264 103420
rect 131264 103400 131266 103420
rect 131394 102720 131450 102776
rect 131118 102176 131174 102232
rect 131210 101088 131266 101144
rect 131210 100408 131266 100464
rect 131118 99864 131174 99920
rect 131210 98640 131266 98696
rect 131118 98096 131174 98152
rect 131210 97552 131266 97608
rect 131670 99320 131726 99376
rect 131578 97008 131634 97064
rect 131210 96328 131266 96384
rect 131118 95784 131174 95840
rect 131394 95240 131450 95296
rect 131210 94560 131266 94616
rect 131118 94016 131174 94072
rect 131210 93472 131266 93528
rect 131118 92792 131174 92848
rect 131210 92248 131266 92304
rect 131118 91704 131174 91760
rect 131210 89936 131266 89992
rect 131210 89392 131266 89448
rect 131118 88712 131174 88768
rect 131210 88204 131212 88224
rect 131212 88204 131264 88224
rect 131264 88204 131266 88224
rect 131210 88168 131266 88204
rect 131118 87624 131174 87680
rect 131302 86944 131358 87000
rect 131118 86400 131174 86456
rect 131210 85856 131266 85912
rect 131210 85312 131266 85368
rect 131118 84632 131174 84688
rect 131210 84108 131266 84144
rect 131210 84088 131212 84108
rect 131212 84088 131264 84108
rect 131264 84088 131266 84108
rect 131578 83544 131634 83600
rect 131118 82864 131174 82920
rect 131210 82320 131266 82376
rect 131118 81776 131174 81832
rect 131210 81096 131266 81152
rect 131118 80552 131174 80608
rect 131210 79908 131212 79928
rect 131212 79908 131264 79928
rect 131264 79908 131266 79928
rect 131210 79872 131266 79908
rect 131118 79464 131174 79520
rect 131302 78784 131358 78840
rect 131210 78240 131266 78296
rect 131118 77696 131174 77752
rect 131210 77052 131212 77072
rect 131212 77052 131264 77072
rect 131264 77052 131266 77072
rect 131210 77016 131266 77052
rect 131302 76472 131358 76528
rect 131670 75928 131726 75984
rect 131210 74704 131266 74760
rect 131210 72936 131266 72992
rect 131118 72392 131174 72448
rect 131302 71848 131358 71904
rect 131210 71168 131266 71224
rect 131118 70624 131174 70680
rect 131210 70080 131266 70136
rect 131118 69400 131174 69456
rect 131210 68892 131212 68912
rect 131212 68892 131264 68912
rect 131264 68892 131266 68912
rect 131210 68856 131266 68892
rect 131394 68312 131450 68368
rect 131118 67768 131174 67824
rect 131210 67088 131266 67144
rect 131118 66544 131174 66600
rect 131210 66000 131266 66056
rect 131118 65320 131174 65376
rect 131210 64796 131266 64832
rect 131210 64776 131212 64796
rect 131212 64776 131264 64796
rect 131264 64776 131266 64796
rect 131302 64232 131358 64288
rect 131118 63688 131174 63744
rect 131210 63008 131266 63064
rect 131210 61956 131212 61976
rect 131212 61956 131264 61976
rect 131264 61956 131266 61976
rect 131210 61920 131266 61956
rect 131118 61240 131174 61296
rect 131210 60152 131266 60208
rect 131118 59472 131174 59528
rect 131578 58928 131634 58984
rect 131210 58384 131266 58440
rect 131210 57876 131212 57896
rect 131212 57876 131264 57896
rect 131264 57876 131266 57896
rect 131210 57840 131266 57876
rect 131210 56616 131266 56672
rect 131210 56072 131266 56128
rect 131118 55392 131174 55448
rect 131210 54304 131266 54360
rect 131210 53660 131212 53680
rect 131212 53660 131264 53680
rect 131264 53660 131266 53680
rect 131210 53624 131266 53660
rect 131670 53080 131726 53136
rect 131118 52536 131174 52592
rect 131210 51312 131266 51368
rect 131210 49544 131266 49600
rect 131302 49000 131358 49056
rect 131210 47232 131266 47288
rect 131118 46144 131174 46200
rect 131210 45484 131266 45520
rect 131210 45464 131212 45484
rect 131212 45464 131264 45484
rect 131264 45464 131266 45484
rect 131118 44376 131174 44432
rect 131210 43696 131266 43752
rect 131210 42644 131212 42664
rect 131212 42644 131264 42664
rect 131264 42644 131266 42664
rect 131210 42608 131266 42644
rect 131118 41928 131174 41984
rect 131210 40840 131266 40896
rect 131118 40296 131174 40352
rect 131210 38564 131212 38584
rect 131212 38564 131264 38584
rect 131264 38564 131266 38584
rect 131210 38528 131266 38564
rect 131118 37848 131174 37904
rect 131670 37304 131726 37360
rect 131302 36760 131358 36816
rect 131210 36080 131266 36136
rect 131210 35536 131266 35592
rect 131118 34992 131174 35048
rect 131210 32680 131266 32736
rect 131118 32000 131174 32056
rect 131210 31456 131266 31512
rect 131302 30912 131358 30968
rect 131118 30368 131174 30424
rect 131946 101632 132002 101688
rect 131854 75248 131910 75304
rect 131854 74160 131910 74216
rect 132314 119720 132370 119776
rect 132314 115640 132370 115696
rect 132222 91160 132278 91216
rect 132222 90480 132278 90536
rect 131946 62464 132002 62520
rect 132038 60696 132094 60752
rect 131854 50224 131910 50280
rect 131946 44920 132002 44976
rect 132314 73616 132370 73672
rect 132222 57160 132278 57216
rect 132130 54848 132186 54904
rect 132222 51992 132278 52048
rect 132130 50768 132186 50824
rect 132314 48456 132370 48512
rect 132038 43152 132094 43208
rect 132222 47776 132278 47832
rect 132406 46688 132462 46744
rect 132130 41384 132186 41440
rect 131854 39616 131910 39672
rect 132498 39072 132554 39128
rect 132130 34448 132186 34504
rect 132038 33768 132094 33824
rect 132222 33224 132278 33280
rect 186318 221176 186374 221232
rect 186318 219952 186374 220008
rect 186318 218864 186374 218920
rect 186410 217776 186466 217832
rect 186318 216708 186374 216744
rect 186318 216688 186320 216708
rect 186320 216688 186372 216708
rect 186372 216688 186374 216708
rect 186318 215464 186374 215520
rect 186318 214376 186374 214432
rect 186318 213288 186374 213344
rect 186318 211148 186320 211168
rect 186320 211148 186372 211168
rect 186372 211148 186374 211168
rect 186318 211112 186374 211148
rect 186318 209888 186374 209944
rect 186318 208664 186374 208720
rect 186318 207576 186374 207632
rect 186318 206488 186374 206544
rect 186318 204332 186374 204368
rect 186318 204312 186320 204332
rect 186320 204312 186372 204332
rect 186372 204312 186374 204332
rect 186318 203088 186374 203144
rect 186318 202000 186374 202056
rect 186318 200776 186374 200832
rect 186410 199688 186466 199744
rect 186318 198756 186374 198792
rect 186318 198736 186320 198756
rect 186320 198736 186372 198756
rect 186372 198736 186374 198756
rect 186318 197512 186374 197568
rect 186318 196288 186374 196344
rect 186318 195200 186374 195256
rect 186318 194112 186374 194168
rect 186410 192888 186466 192944
rect 186318 191836 186320 191856
rect 186320 191836 186372 191856
rect 186372 191836 186374 191856
rect 186318 191800 186374 191836
rect 186318 190712 186374 190768
rect 186318 189488 186374 189544
rect 186318 188400 186374 188456
rect 186410 187312 186466 187368
rect 186318 186396 186320 186416
rect 186320 186396 186372 186416
rect 186372 186396 186374 186416
rect 186318 186360 186374 186396
rect 186318 183912 186374 183968
rect 186318 182824 186374 182880
rect 186318 181600 186374 181656
rect 186410 180512 186466 180568
rect 186318 179460 186320 179480
rect 186320 179460 186372 179480
rect 186372 179460 186374 179480
rect 186318 179424 186374 179460
rect 186318 178200 186374 178256
rect 186318 177112 186374 177168
rect 186318 176024 186374 176080
rect 186318 174936 186374 174992
rect 186318 172624 186374 172680
rect 186318 171536 186374 171592
rect 186318 170312 186374 170368
rect 186318 169224 186374 169280
rect 186410 168136 186466 168192
rect 186318 167084 186320 167104
rect 186320 167084 186372 167104
rect 186372 167084 186374 167104
rect 186318 167048 186374 167084
rect 186318 165824 186374 165880
rect 186318 164736 186374 164792
rect 186318 163648 186374 163704
rect 186410 162424 186466 162480
rect 186318 161508 186320 161528
rect 186320 161508 186372 161528
rect 186372 161508 186374 161528
rect 186318 161472 186374 161508
rect 186318 160248 186374 160304
rect 186318 159024 186374 159080
rect 186318 157936 186374 157992
rect 186318 156848 186374 156904
rect 186410 155760 186466 155816
rect 186318 154692 186374 154728
rect 186318 154672 186320 154692
rect 186320 154672 186372 154692
rect 186372 154672 186374 154692
rect 186318 153448 186374 153504
rect 186318 152360 186374 152416
rect 186318 151136 186374 151192
rect 186410 150048 186466 150104
rect 186318 149132 186320 149152
rect 186320 149132 186372 149152
rect 186372 149132 186374 149152
rect 186318 149096 186374 149132
rect 186318 147736 186374 147792
rect 186318 146648 186374 146704
rect 186318 145560 186374 145616
rect 186318 144472 186374 144528
rect 186410 143248 186466 143304
rect 186318 142180 186374 142216
rect 186318 142160 186320 142180
rect 186320 142160 186372 142180
rect 186372 142160 186374 142180
rect 186318 139848 186374 139904
rect 186318 138760 186374 138816
rect 186318 137672 186374 137728
rect 186410 136448 186466 136504
rect 186318 135380 186374 135416
rect 186318 135360 186320 135380
rect 186320 135360 186372 135380
rect 186372 135360 186374 135380
rect 186318 134272 186374 134328
rect 186318 133184 186374 133240
rect 186318 131960 186374 132016
rect 133142 28872 133198 28928
rect 131762 28736 131818 28792
rect 186318 129804 186374 129840
rect 186318 129784 186320 129804
rect 186320 129784 186372 129804
rect 186372 129784 186374 129804
rect 186318 128560 186374 128616
rect 186318 127472 186374 127528
rect 186318 126384 186374 126440
rect 186318 125160 186374 125216
rect 186318 122984 186374 123040
rect 186318 121896 186374 121952
rect 186318 119584 186374 119640
rect 186410 118496 186466 118552
rect 186318 117308 186320 117328
rect 186320 117308 186372 117328
rect 186372 117308 186374 117328
rect 186318 117272 186374 117308
rect 186318 116184 186374 116240
rect 186318 115096 186374 115152
rect 186318 114008 186374 114064
rect 186410 112784 186466 112840
rect 186318 111852 186374 111888
rect 186318 111832 186320 111852
rect 186320 111832 186372 111852
rect 186372 111832 186374 111852
rect 186318 109384 186374 109440
rect 186318 108296 186374 108352
rect 186318 107208 186374 107264
rect 186410 105984 186466 106040
rect 186318 104916 186374 104952
rect 186318 104896 186320 104916
rect 186320 104896 186372 104916
rect 186372 104896 186374 104916
rect 186318 102720 186374 102776
rect 186318 101496 186374 101552
rect 186410 100408 186466 100464
rect 186318 99456 186374 99512
rect 186318 98096 186374 98152
rect 186318 97008 186374 97064
rect 186318 95920 186374 95976
rect 186318 94696 186374 94752
rect 186410 93608 186466 93664
rect 186318 92540 186374 92576
rect 186318 92520 186320 92540
rect 186320 92520 186372 92540
rect 186372 92520 186374 92540
rect 186318 91432 186374 91488
rect 186318 90208 186374 90264
rect 186318 89120 186374 89176
rect 186318 88032 186374 88088
rect 186318 85720 186374 85776
rect 186318 84632 186374 84688
rect 186318 82320 186374 82376
rect 186318 81232 186374 81288
rect 186318 78920 186374 78976
rect 186318 77832 186374 77888
rect 186410 75520 186466 75576
rect 186318 74588 186374 74624
rect 186318 74568 186320 74588
rect 186320 74568 186372 74588
rect 186372 74568 186374 74588
rect 186318 72256 186374 72312
rect 186318 71032 186374 71088
rect 186318 69944 186374 70000
rect 186410 69028 186412 69048
rect 186412 69028 186464 69048
rect 186464 69028 186466 69048
rect 186410 68992 186466 69028
rect 186318 67652 186374 67688
rect 186318 67632 186320 67652
rect 186320 67632 186372 67652
rect 186372 67632 186374 67652
rect 186318 66544 186374 66600
rect 186318 65456 186374 65512
rect 186318 64232 186374 64288
rect 186318 62192 186374 62248
rect 186318 60968 186374 61024
rect 186318 58656 186374 58712
rect 186318 57568 186374 57624
rect 186318 55276 186374 55312
rect 186318 55256 186320 55276
rect 186320 55256 186372 55276
rect 186372 55256 186374 55276
rect 186318 54168 186374 54224
rect 186318 51856 186374 51912
rect 186318 50768 186374 50824
rect 186318 48456 186374 48512
rect 186318 47368 186374 47424
rect 186594 45056 186650 45112
rect 186410 43968 186466 44024
rect 186318 42880 186374 42936
rect 186502 41656 186558 41712
rect 186410 38392 186466 38448
rect 186318 37324 186374 37360
rect 186318 37304 186320 37324
rect 186320 37304 186372 37324
rect 186372 37304 186374 37324
rect 186318 36080 186374 36136
rect 186410 34992 186466 35048
rect 186318 33768 186374 33824
rect 186410 32680 186466 32736
rect 186318 31728 186374 31784
rect 186318 30504 186374 30560
rect 187514 224712 187570 224768
rect 187606 223488 187662 223544
rect 186962 212064 187018 212120
rect 187054 205400 187110 205456
rect 187146 185000 187202 185056
rect 186962 120672 187018 120728
rect 187054 110608 187110 110664
rect 186962 73344 187018 73400
rect 187238 173712 187294 173768
rect 187330 141072 187386 141128
rect 187146 103808 187202 103864
rect 187422 130872 187478 130928
rect 187238 86944 187294 87000
rect 187146 63144 187202 63200
rect 187054 59744 187110 59800
rect 186962 49680 187018 49736
rect 187330 83408 187386 83464
rect 187514 124208 187570 124264
rect 187422 80144 187478 80200
rect 187514 76744 187570 76800
rect 187238 56344 187294 56400
rect 187146 46280 187202 46336
rect 186962 39480 187018 39536
rect 187330 52944 187386 53000
rect 187238 40568 187294 40624
rect 207018 307128 207074 307184
rect 207018 305496 207074 305552
rect 209686 332832 209742 332888
rect 209594 331064 209650 331120
rect 238666 299784 238722 299840
rect 215850 298016 215906 298072
rect 224958 298016 225014 298072
rect 226338 298016 226394 298072
rect 227718 298016 227774 298072
rect 229190 298016 229246 298072
rect 230478 298016 230534 298072
rect 231858 298016 231914 298072
rect 233238 298016 233294 298072
rect 234618 298016 234674 298072
rect 237194 298016 237250 298072
rect 229466 297200 229522 297256
rect 237378 297880 237434 297936
rect 237286 297744 237342 297800
rect 243082 299648 243138 299704
rect 238758 298016 238814 298072
rect 240138 298016 240194 298072
rect 241426 298016 241482 298072
rect 242898 298016 242954 298072
rect 238666 297064 238722 297120
rect 238666 296792 238722 296848
rect 240046 297064 240102 297120
rect 241518 297880 241574 297936
rect 242806 297744 242862 297800
rect 244094 298016 244150 298072
rect 244278 298016 244334 298072
rect 245566 298016 245622 298072
rect 246854 298016 246910 298072
rect 248326 298016 248382 298072
rect 249706 298016 249762 298072
rect 251086 298016 251142 298072
rect 252374 298016 252430 298072
rect 253754 298016 253810 298072
rect 255134 298016 255190 298072
rect 256514 298016 256570 298072
rect 257802 298016 257858 298072
rect 257986 298016 258042 298072
rect 259182 298016 259238 298072
rect 260654 298016 260710 298072
rect 262034 298016 262090 298072
rect 263506 298016 263562 298072
rect 266174 298016 266230 298072
rect 273166 298016 273222 298072
rect 274546 298016 274602 298072
rect 275926 298016 275982 298072
rect 277306 298016 277362 298072
rect 243082 297880 243138 297936
rect 244186 297880 244242 297936
rect 246762 297880 246818 297936
rect 248234 297880 248290 297936
rect 246946 297744 247002 297800
rect 249614 297880 249670 297936
rect 250994 297880 251050 297936
rect 252282 297880 252338 297936
rect 252466 297744 252522 297800
rect 253846 297880 253902 297936
rect 255226 297880 255282 297936
rect 256606 297880 256662 297936
rect 257894 297880 257950 297936
rect 259366 297880 259422 297936
rect 259274 297744 259330 297800
rect 260746 297880 260802 297936
rect 262126 297880 262182 297936
rect 263414 297880 263470 297936
rect 264794 296928 264850 296984
rect 264886 296792 264942 296848
rect 269026 297472 269082 297528
rect 267554 297064 267610 297120
rect 266266 296792 266322 296848
rect 267462 296792 267518 296848
rect 267646 296928 267702 296984
rect 270406 296792 270462 296848
rect 271786 296792 271842 296848
rect 273074 296792 273130 296848
rect 408498 249600 408554 249656
rect 409326 247696 409382 247752
rect 409326 233688 409382 233744
rect 409326 231784 409382 231840
rect 409326 230016 409382 230072
rect 410062 226072 410118 226128
rect 409970 223216 410026 223272
rect 411258 245112 411314 245168
rect 410522 243208 410578 243264
rect 410430 241168 410486 241224
rect 411258 235320 411314 235376
rect 410338 227432 410394 227488
rect 410246 221584 410302 221640
rect 410154 217640 410210 217696
rect 411626 239264 411682 239320
rect 411534 237224 411590 237280
rect 579618 232328 579674 232384
rect 411718 219544 411774 219600
rect 411442 215600 411498 215656
rect 411350 213696 411406 213752
rect 409878 212336 409934 212392
rect 411258 209788 411260 209808
rect 411260 209788 411312 209808
rect 411312 209788 411314 209808
rect 411258 209752 411314 209788
rect 411258 207848 411314 207904
rect 411258 205808 411314 205864
rect 411258 203904 411314 203960
rect 411902 201864 411958 201920
rect 411258 197920 411314 197976
rect 411258 196036 411314 196072
rect 411258 196016 411260 196036
rect 411260 196016 411312 196036
rect 411312 196016 411314 196036
rect 411258 192072 411314 192128
rect 411258 190168 411314 190224
rect 411258 188128 411314 188184
rect 411258 186224 411314 186280
rect 411258 184184 411314 184240
rect 411258 182280 411314 182336
rect 411258 180240 411314 180296
rect 411258 178336 411314 178392
rect 411258 176432 411314 176488
rect 411258 174392 411314 174448
rect 411258 172524 411260 172544
rect 411260 172524 411312 172544
rect 411312 172524 411314 172544
rect 411258 172488 411314 172524
rect 411258 170448 411314 170504
rect 411258 168544 411314 168600
rect 411258 166504 411314 166560
rect 411258 164600 411314 164656
rect 411258 162560 411314 162616
rect 411258 160656 411314 160712
rect 411258 158772 411314 158808
rect 411258 158752 411260 158772
rect 411260 158752 411312 158772
rect 411312 158752 411314 158772
rect 411258 156712 411314 156768
rect 411258 154808 411314 154864
rect 411258 152768 411314 152824
rect 411258 150864 411314 150920
rect 411258 148824 411314 148880
rect 411258 146920 411314 146976
rect 411258 144916 411260 144936
rect 411260 144916 411312 144936
rect 411312 144916 411314 144936
rect 411258 144880 411314 144916
rect 411258 142976 411314 143032
rect 411258 141072 411314 141128
rect 411258 139032 411314 139088
rect 411258 137128 411314 137184
rect 411258 135088 411314 135144
rect 411258 133184 411314 133240
rect 411258 129240 411314 129296
rect 411258 127200 411314 127256
rect 411258 125296 411314 125352
rect 411258 123256 411314 123312
rect 411258 121352 411314 121408
rect 411258 119448 411314 119504
rect 411258 115504 411314 115560
rect 412086 199960 412142 200016
rect 411994 194112 412050 194168
rect 411258 113464 411314 113520
rect 411902 111560 411958 111616
rect 411258 109520 411314 109576
rect 411258 107652 411260 107672
rect 411260 107652 411312 107672
rect 411312 107652 411314 107672
rect 411258 107616 411314 107652
rect 411258 103672 411314 103728
rect 411258 101768 411314 101824
rect 411258 95820 411260 95840
rect 411260 95820 411312 95840
rect 411312 95820 411314 95840
rect 411258 95784 411314 95820
rect 411258 93916 411260 93936
rect 411260 93916 411312 93936
rect 411312 93916 411314 93936
rect 411258 93880 411314 93916
rect 411258 91840 411314 91896
rect 411258 89936 411314 89992
rect 411258 87896 411314 87952
rect 411258 85992 411314 86048
rect 411258 84124 411260 84144
rect 411260 84124 411312 84144
rect 411312 84124 411314 84144
rect 411258 84088 411314 84124
rect 411258 82048 411314 82104
rect 411258 78104 411314 78160
rect 411258 76200 411314 76256
rect 411258 74196 411260 74216
rect 411260 74196 411312 74216
rect 411312 74196 411314 74216
rect 411258 74160 411314 74196
rect 411258 72256 411314 72312
rect 411350 70216 411406 70272
rect 411258 68312 411314 68368
rect 411258 66408 411314 66464
rect 411258 64368 411314 64424
rect 411258 62464 411314 62520
rect 411258 60424 411314 60480
rect 411258 58520 411314 58576
rect 411258 54576 411314 54632
rect 411258 52556 411314 52592
rect 411258 52536 411260 52556
rect 411260 52536 411312 52556
rect 411312 52536 411314 52556
rect 411258 48728 411314 48784
rect 411258 42744 411314 42800
rect 412178 131144 412234 131200
rect 411994 105576 412050 105632
rect 411258 40840 411314 40896
rect 411258 38836 411260 38856
rect 411260 38836 411312 38856
rect 411312 38836 411314 38856
rect 411258 38800 411314 38836
rect 411258 36896 411314 36952
rect 411258 34856 411314 34912
rect 411258 32952 411314 33008
rect 411258 31048 411314 31104
rect 412086 99728 412142 99784
rect 412270 117408 412326 117464
rect 412178 56480 412234 56536
rect 412362 97824 412418 97880
rect 412270 44784 412326 44840
rect 412546 80144 412602 80200
rect 412454 50632 412510 50688
rect 412546 46688 412602 46744
rect 405738 28872 405794 28928
rect 397458 28736 397514 28792
rect 580170 219000 580226 219056
rect 437478 128696 437534 128752
rect 437478 127336 437534 127392
rect 539322 125976 539378 126032
rect 437478 125840 437534 125896
rect 437478 124228 437534 124264
rect 437478 124208 437480 124228
rect 437480 124208 437532 124228
rect 437532 124208 437534 124228
rect 437478 122984 437534 123040
rect 438490 120808 438546 120864
rect 436742 106120 436798 106176
rect 438398 119176 438454 119232
rect 438306 117680 438362 117736
rect 438214 116048 438270 116104
rect 438122 114552 438178 114608
rect 437478 114008 437534 114064
rect 437478 112512 437534 112568
rect 437478 110200 437534 110256
rect 437478 108996 437534 109032
rect 437478 108976 437480 108996
rect 437480 108976 437532 108996
rect 437532 108976 437534 108996
rect 437478 107344 437534 107400
rect 437478 104488 437534 104544
rect 437662 103028 437664 103048
rect 437664 103028 437716 103048
rect 437716 103028 437718 103048
rect 437662 102992 437718 103028
rect 437478 101496 437534 101552
rect 437478 100000 437534 100056
rect 437478 97688 437534 97744
rect 437478 96464 437534 96520
rect 437478 95140 437480 95160
rect 437480 95140 437532 95160
rect 437532 95140 437534 95160
rect 437478 95104 437534 95140
rect 437478 93472 437534 93528
rect 437478 91976 437534 92032
rect 437478 90480 437534 90536
rect 437478 88984 437534 89040
rect 437478 87488 437534 87544
rect 437478 85484 437480 85504
rect 437480 85484 437532 85504
rect 437532 85484 437534 85504
rect 437478 85448 437534 85484
rect 437478 84124 437480 84144
rect 437480 84124 437532 84144
rect 437532 84124 437534 84144
rect 437478 84088 437534 84124
rect 437478 82456 437534 82512
rect 437478 80960 437534 81016
rect 437478 79600 437534 79656
rect 437478 78104 437534 78160
rect 437478 76608 437534 76664
rect 437478 74296 437534 74352
rect 437478 73092 437534 73128
rect 437478 73072 437480 73092
rect 437480 73072 437532 73092
rect 437532 73072 437534 73092
rect 437478 71440 437534 71496
rect 437478 70216 437534 70272
rect 437478 68584 437534 68640
rect 437478 67088 437534 67144
rect 437478 65592 437534 65648
rect 437478 64096 437534 64152
rect 437478 62076 437534 62112
rect 437478 62056 437480 62076
rect 437480 62056 437532 62076
rect 437532 62056 437534 62076
rect 437478 60560 437534 60616
rect 437478 59200 437534 59256
rect 437478 57568 437534 57624
rect 437478 56072 437534 56128
rect 437754 54576 437810 54632
rect 437478 53080 437534 53136
rect 437478 51584 437534 51640
rect 436834 49544 436890 49600
rect 437478 48220 437480 48240
rect 437480 48220 437532 48240
rect 437532 48220 437534 48240
rect 437478 48184 437534 48220
rect 437478 46552 437534 46608
rect 437478 45192 437534 45248
rect 437478 43560 437534 43616
rect 437478 42200 437534 42256
rect 437478 40568 437534 40624
rect 437478 38392 437534 38448
rect 437478 37204 437480 37224
rect 437480 37204 437532 37224
rect 437532 37204 437534 37224
rect 437478 37168 437534 37204
rect 437478 35844 437480 35864
rect 437480 35844 437532 35864
rect 437532 35844 437534 35864
rect 437478 35808 437534 35844
rect 437478 34040 437534 34096
rect 542450 116320 542506 116376
rect 542358 107208 542414 107264
rect 542358 98096 542414 98152
rect 437478 32680 437534 32736
rect 437478 31184 437534 31240
rect 542450 88984 542506 89040
rect 542542 80008 542598 80064
rect 542634 70896 542690 70952
rect 542726 61784 542782 61840
rect 543002 43560 543058 43616
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580354 152632 580410 152688
rect 580354 125976 580410 126032
rect 580262 112784 580318 112840
rect 580170 99456 580226 99512
rect 580262 86128 580318 86184
rect 579802 59608 579858 59664
rect 543186 52672 543242 52728
rect 543094 34584 543150 34640
rect 580170 33088 580226 33144
rect 580446 72936 580502 72992
rect 580538 46280 580594 46336
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect 48221 334250 48287 334253
rect 48221 334248 49434 334250
rect 48221 334192 48226 334248
rect 48282 334204 49434 334248
rect 48282 334192 50048 334204
rect 48221 334190 50048 334192
rect 48221 334187 48287 334190
rect 49374 334144 50048 334190
rect 209730 334144 210032 334204
rect 208301 334114 208367 334117
rect 209730 334114 209790 334144
rect 208301 334112 209790 334114
rect 208301 334056 208306 334112
rect 208362 334056 209790 334112
rect 208301 334054 209790 334056
rect 208301 334051 208367 334054
rect 48129 333026 48195 333029
rect 48129 333024 49434 333026
rect 48129 332968 48134 333024
rect 48190 332980 49434 333024
rect 48190 332968 50048 332980
rect 48129 332966 50048 332968
rect 48129 332963 48195 332966
rect 49374 332920 50048 332966
rect 209730 332920 210032 332980
rect 209730 332893 209790 332920
rect 209681 332888 209790 332893
rect 209681 332832 209686 332888
rect 209742 332832 209790 332888
rect 209681 332830 209790 332832
rect 209681 332827 209747 332830
rect -960 332196 480 332436
rect 49742 331152 50048 331212
rect 209730 331152 210032 331212
rect 47945 331122 48011 331125
rect 49742 331122 49802 331152
rect 47945 331120 49802 331122
rect 47945 331064 47950 331120
rect 48006 331064 49802 331120
rect 47945 331062 49802 331064
rect 209589 331122 209655 331125
rect 209730 331122 209790 331152
rect 209589 331120 209790 331122
rect 209589 331064 209594 331120
rect 209650 331064 209790 331120
rect 209589 331062 209790 331064
rect 47945 331059 48011 331062
rect 209589 331059 209655 331062
rect 49601 330124 49667 330127
rect 49601 330122 50048 330124
rect 49601 330066 49606 330122
rect 49662 330066 50048 330122
rect 49601 330064 50048 330066
rect 209730 330064 210032 330124
rect 49601 330061 49667 330064
rect 208209 330034 208275 330037
rect 209730 330034 209790 330064
rect 208209 330032 209790 330034
rect 208209 329976 208214 330032
rect 208270 329976 209790 330032
rect 208209 329974 209790 329976
rect 208209 329971 208275 329974
rect 47853 328538 47919 328541
rect 208117 328538 208183 328541
rect 47853 328536 49434 328538
rect 47853 328480 47858 328536
rect 47914 328492 49434 328536
rect 208117 328536 209790 328538
rect 47914 328480 50048 328492
rect 47853 328478 50048 328480
rect 47853 328475 47919 328478
rect 49374 328432 50048 328478
rect 208117 328480 208122 328536
rect 208178 328492 209790 328536
rect 208178 328480 210032 328492
rect 208117 328478 210032 328480
rect 208117 328475 208183 328478
rect 209730 328432 210032 328478
rect 47761 327586 47827 327589
rect 47761 327584 49434 327586
rect 47761 327528 47766 327584
rect 47822 327540 49434 327584
rect 47822 327528 50048 327540
rect 47761 327526 50048 327528
rect 47761 327523 47827 327526
rect 49374 327480 50048 327526
rect 209730 327480 210032 327540
rect 208025 327450 208091 327453
rect 209730 327450 209790 327480
rect 208025 327448 209790 327450
rect 208025 327392 208030 327448
rect 208086 327392 209790 327448
rect 208025 327390 209790 327392
rect 208025 327387 208091 327390
rect 48037 325818 48103 325821
rect 207013 325818 207079 325821
rect 48037 325816 49434 325818
rect 48037 325760 48042 325816
rect 48098 325772 49434 325816
rect 207013 325816 209790 325818
rect 48098 325760 50048 325772
rect 48037 325758 50048 325760
rect 48037 325755 48103 325758
rect 49374 325712 50048 325758
rect 207013 325760 207018 325816
rect 207074 325772 209790 325816
rect 207074 325760 210032 325772
rect 207013 325758 210032 325760
rect 207013 325755 207079 325758
rect 209730 325712 210032 325758
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect 49509 307276 49575 307279
rect 49509 307274 50048 307276
rect 49509 307218 49514 307274
rect 49570 307218 50048 307274
rect 49509 307216 50048 307218
rect 209730 307216 210032 307276
rect 49509 307213 49575 307216
rect 207013 307186 207079 307189
rect 209730 307186 209790 307216
rect 207013 307184 209790 307186
rect 207013 307128 207018 307184
rect 207074 307128 209790 307184
rect 207013 307126 209790 307128
rect 207013 307123 207079 307126
rect -960 306084 480 306324
rect 47669 305690 47735 305693
rect 47669 305688 49434 305690
rect 47669 305632 47674 305688
rect 47730 305644 49434 305688
rect 47730 305632 50048 305644
rect 47669 305630 50048 305632
rect 47669 305627 47735 305630
rect 49374 305584 50048 305630
rect 209730 305584 210032 305644
rect 207013 305554 207079 305557
rect 209730 305554 209790 305584
rect 207013 305552 209790 305554
rect 207013 305496 207018 305552
rect 207074 305496 209790 305552
rect 207013 305494 209790 305496
rect 207013 305491 207079 305494
rect 238661 299842 238727 299845
rect 239648 299842 239654 299844
rect 238661 299840 239654 299842
rect 238661 299784 238666 299840
rect 238722 299784 239654 299840
rect 238661 299782 239654 299784
rect 238661 299779 238727 299782
rect 239648 299780 239654 299782
rect 239718 299780 239724 299844
rect 243077 299708 243143 299709
rect 243048 299706 243054 299708
rect 242986 299646 243054 299706
rect 243118 299704 243143 299708
rect 243138 299648 243143 299704
rect 243048 299644 243054 299646
rect 243118 299644 243143 299648
rect 243077 299643 243143 299644
rect 55857 299572 55923 299573
rect 55848 299570 55854 299572
rect 55766 299510 55854 299570
rect 55848 299508 55854 299510
rect 55918 299508 55924 299572
rect 55857 299507 55923 299508
rect 583520 298604 584960 298844
rect 103237 298212 103303 298213
rect 73654 298148 73660 298212
rect 73724 298148 73730 298212
rect 77886 298148 77892 298212
rect 77956 298148 77962 298212
rect 81750 298148 81756 298212
rect 81820 298148 81826 298212
rect 85430 298148 85436 298212
rect 85500 298148 85506 298212
rect 91870 298148 91876 298212
rect 91940 298148 91946 298212
rect 95550 298148 95556 298212
rect 95620 298148 95626 298212
rect 95918 298148 95924 298212
rect 95988 298148 95994 298212
rect 99414 298148 99420 298212
rect 99484 298148 99490 298212
rect 102910 298148 102916 298212
rect 102980 298148 102986 298212
rect 103237 298208 103284 298212
rect 103348 298210 103354 298212
rect 103237 298152 103242 298208
rect 103237 298148 103284 298152
rect 103348 298150 103394 298210
rect 103348 298148 103354 298150
rect 225454 298148 225460 298212
rect 225524 298148 225530 298212
rect 229134 298148 229140 298212
rect 229204 298148 229210 298212
rect 257838 298148 257844 298212
rect 257908 298210 257914 298212
rect 257908 298150 258090 298210
rect 257908 298148 257914 298150
rect 65558 298012 65564 298076
rect 65628 298074 65634 298076
rect 65701 298074 65767 298077
rect 65628 298072 65767 298074
rect 65628 298016 65706 298072
rect 65762 298016 65767 298072
rect 65628 298014 65767 298016
rect 65628 298012 65634 298014
rect 65701 298011 65767 298014
rect 66662 298012 66668 298076
rect 66732 298074 66738 298076
rect 67541 298074 67607 298077
rect 67817 298076 67883 298077
rect 66732 298072 67607 298074
rect 66732 298016 67546 298072
rect 67602 298016 67607 298072
rect 66732 298014 67607 298016
rect 66732 298012 66738 298014
rect 67541 298011 67607 298014
rect 67766 298012 67772 298076
rect 67836 298074 67883 298076
rect 67836 298072 67928 298074
rect 67878 298016 67928 298072
rect 67836 298014 67928 298016
rect 67836 298012 67883 298014
rect 69238 298012 69244 298076
rect 69308 298074 69314 298076
rect 69933 298074 69999 298077
rect 70209 298076 70275 298077
rect 71497 298076 71563 298077
rect 70158 298074 70164 298076
rect 69308 298072 69999 298074
rect 69308 298016 69938 298072
rect 69994 298016 69999 298072
rect 69308 298014 69999 298016
rect 70118 298014 70164 298074
rect 70228 298072 70275 298076
rect 71446 298074 71452 298076
rect 70270 298016 70275 298072
rect 69308 298012 69314 298014
rect 67817 298011 67883 298012
rect 69933 298011 69999 298014
rect 70158 298012 70164 298014
rect 70228 298012 70275 298016
rect 71406 298014 71452 298074
rect 71516 298072 71563 298076
rect 71558 298016 71563 298072
rect 71446 298012 71452 298014
rect 71516 298012 71563 298016
rect 72550 298012 72556 298076
rect 72620 298074 72626 298076
rect 73061 298074 73127 298077
rect 72620 298072 73127 298074
rect 72620 298016 73066 298072
rect 73122 298016 73127 298072
rect 72620 298014 73127 298016
rect 73662 298074 73722 298148
rect 74441 298074 74507 298077
rect 73662 298072 74507 298074
rect 73662 298016 74446 298072
rect 74502 298016 74507 298072
rect 73662 298014 74507 298016
rect 72620 298012 72626 298014
rect 70209 298011 70275 298012
rect 71497 298011 71563 298012
rect 73061 298011 73127 298014
rect 74441 298011 74507 298014
rect 75126 298012 75132 298076
rect 75196 298074 75202 298076
rect 75821 298074 75887 298077
rect 75196 298072 75887 298074
rect 75196 298016 75826 298072
rect 75882 298016 75887 298072
rect 75196 298014 75887 298016
rect 75196 298012 75202 298014
rect 75821 298011 75887 298014
rect 76230 298012 76236 298076
rect 76300 298074 76306 298076
rect 76833 298074 76899 298077
rect 76300 298072 76899 298074
rect 76300 298016 76838 298072
rect 76894 298016 76899 298072
rect 76300 298014 76899 298016
rect 76300 298012 76306 298014
rect 76833 298011 76899 298014
rect 77109 298076 77175 298077
rect 77109 298072 77156 298076
rect 77220 298074 77226 298076
rect 77109 298016 77114 298072
rect 77109 298012 77156 298016
rect 77220 298014 77266 298074
rect 77220 298012 77226 298014
rect 77109 298011 77175 298012
rect 77894 297938 77954 298148
rect 81758 298077 81818 298148
rect 78254 298012 78260 298076
rect 78324 298074 78330 298076
rect 78581 298074 78647 298077
rect 78324 298072 78647 298074
rect 78324 298016 78586 298072
rect 78642 298016 78647 298072
rect 78324 298014 78647 298016
rect 78324 298012 78330 298014
rect 78581 298011 78647 298014
rect 79358 298012 79364 298076
rect 79428 298074 79434 298076
rect 79869 298074 79935 298077
rect 79428 298072 79935 298074
rect 79428 298016 79874 298072
rect 79930 298016 79935 298072
rect 79428 298014 79935 298016
rect 79428 298012 79434 298014
rect 79869 298011 79935 298014
rect 80830 298012 80836 298076
rect 80900 298074 80906 298076
rect 81249 298074 81315 298077
rect 80900 298072 81315 298074
rect 80900 298016 81254 298072
rect 81310 298016 81315 298072
rect 80900 298014 81315 298016
rect 81758 298072 81867 298077
rect 81758 298016 81806 298072
rect 81862 298016 81867 298072
rect 81758 298014 81867 298016
rect 80900 298012 80906 298014
rect 81249 298011 81315 298014
rect 81801 298011 81867 298014
rect 82118 298012 82124 298076
rect 82188 298074 82194 298076
rect 82629 298074 82695 298077
rect 82188 298072 82695 298074
rect 82188 298016 82634 298072
rect 82690 298016 82695 298072
rect 82188 298014 82695 298016
rect 82188 298012 82194 298014
rect 82629 298011 82695 298014
rect 83222 298012 83228 298076
rect 83292 298074 83298 298076
rect 84009 298074 84075 298077
rect 83292 298072 84075 298074
rect 83292 298016 84014 298072
rect 84070 298016 84075 298072
rect 83292 298014 84075 298016
rect 83292 298012 83298 298014
rect 84009 298011 84075 298014
rect 84510 298012 84516 298076
rect 84580 298074 84586 298076
rect 85297 298074 85363 298077
rect 84580 298072 85363 298074
rect 84580 298016 85302 298072
rect 85358 298016 85363 298072
rect 84580 298014 85363 298016
rect 84580 298012 84586 298014
rect 85297 298011 85363 298014
rect 85438 297941 85498 298148
rect 86534 298012 86540 298076
rect 86604 298074 86610 298076
rect 86769 298074 86835 298077
rect 86604 298072 86835 298074
rect 86604 298016 86774 298072
rect 86830 298016 86835 298072
rect 86604 298014 86835 298016
rect 86604 298012 86610 298014
rect 86769 298011 86835 298014
rect 87822 298012 87828 298076
rect 87892 298074 87898 298076
rect 88149 298074 88215 298077
rect 87892 298072 88215 298074
rect 87892 298016 88154 298072
rect 88210 298016 88215 298072
rect 87892 298014 88215 298016
rect 87892 298012 87898 298014
rect 88149 298011 88215 298014
rect 89294 298012 89300 298076
rect 89364 298074 89370 298076
rect 89621 298074 89687 298077
rect 89364 298072 89687 298074
rect 89364 298016 89626 298072
rect 89682 298016 89687 298072
rect 89364 298014 89687 298016
rect 89364 298012 89370 298014
rect 89621 298011 89687 298014
rect 90766 298012 90772 298076
rect 90836 298074 90842 298076
rect 90909 298074 90975 298077
rect 90836 298072 90975 298074
rect 90836 298016 90914 298072
rect 90970 298016 90975 298072
rect 90836 298014 90975 298016
rect 91878 298074 91938 298148
rect 92381 298074 92447 298077
rect 91878 298072 92447 298074
rect 91878 298016 92386 298072
rect 92442 298016 92447 298072
rect 91878 298014 92447 298016
rect 90836 298012 90842 298014
rect 90909 298011 90975 298014
rect 92381 298011 92447 298014
rect 93158 298012 93164 298076
rect 93228 298074 93234 298076
rect 93301 298074 93367 298077
rect 93228 298072 93367 298074
rect 93228 298016 93306 298072
rect 93362 298016 93367 298072
rect 93228 298014 93367 298016
rect 93228 298012 93234 298014
rect 93301 298011 93367 298014
rect 93526 298012 93532 298076
rect 93596 298074 93602 298076
rect 93669 298074 93735 298077
rect 93596 298072 93735 298074
rect 93596 298016 93674 298072
rect 93730 298016 93735 298072
rect 93596 298014 93735 298016
rect 93596 298012 93602 298014
rect 93669 298011 93735 298014
rect 94446 298012 94452 298076
rect 94516 298074 94522 298076
rect 95049 298074 95115 298077
rect 94516 298072 95115 298074
rect 94516 298016 95054 298072
rect 95110 298016 95115 298072
rect 94516 298014 95115 298016
rect 94516 298012 94522 298014
rect 95049 298011 95115 298014
rect 78489 297938 78555 297941
rect 79777 297940 79843 297941
rect 79726 297938 79732 297940
rect 77894 297936 78555 297938
rect 77894 297880 78494 297936
rect 78550 297880 78555 297936
rect 77894 297878 78555 297880
rect 79686 297878 79732 297938
rect 79796 297936 79843 297940
rect 79838 297880 79843 297936
rect 78489 297875 78555 297878
rect 79726 297876 79732 297878
rect 79796 297876 79843 297880
rect 80278 297876 80284 297940
rect 80348 297938 80354 297940
rect 81341 297938 81407 297941
rect 80348 297936 81407 297938
rect 80348 297880 81346 297936
rect 81402 297880 81407 297936
rect 80348 297878 81407 297880
rect 80348 297876 80354 297878
rect 79777 297875 79843 297876
rect 81341 297875 81407 297878
rect 83038 297876 83044 297940
rect 83108 297938 83114 297940
rect 84101 297938 84167 297941
rect 83108 297936 84167 297938
rect 83108 297880 84106 297936
rect 84162 297880 84167 297936
rect 83108 297878 84167 297880
rect 83108 297876 83114 297878
rect 84101 297875 84167 297878
rect 85389 297936 85498 297941
rect 85389 297880 85394 297936
rect 85450 297880 85498 297936
rect 85389 297878 85498 297880
rect 86677 297938 86743 297941
rect 86902 297938 86908 297940
rect 86677 297936 86908 297938
rect 86677 297880 86682 297936
rect 86738 297880 86908 297936
rect 86677 297878 86908 297880
rect 85389 297875 85455 297878
rect 86677 297875 86743 297878
rect 86902 297876 86908 297878
rect 86972 297876 86978 297940
rect 87638 297876 87644 297940
rect 87708 297938 87714 297940
rect 88241 297938 88307 297941
rect 87708 297936 88307 297938
rect 87708 297880 88246 297936
rect 88302 297880 88307 297936
rect 87708 297878 88307 297880
rect 87708 297876 87714 297878
rect 88241 297875 88307 297878
rect 88926 297876 88932 297940
rect 88996 297938 89002 297940
rect 89529 297938 89595 297941
rect 88996 297936 89595 297938
rect 88996 297880 89534 297936
rect 89590 297880 89595 297936
rect 88996 297878 89595 297880
rect 88996 297876 89002 297878
rect 89529 297875 89595 297878
rect 90214 297876 90220 297940
rect 90284 297938 90290 297940
rect 91001 297938 91067 297941
rect 90284 297936 91067 297938
rect 90284 297880 91006 297936
rect 91062 297880 91067 297936
rect 90284 297878 91067 297880
rect 90284 297876 90290 297878
rect 91001 297875 91067 297878
rect 91318 297876 91324 297940
rect 91388 297938 91394 297940
rect 92289 297938 92355 297941
rect 91388 297936 92355 297938
rect 91388 297880 92294 297936
rect 92350 297880 92355 297936
rect 91388 297878 92355 297880
rect 91388 297876 91394 297878
rect 92289 297875 92355 297878
rect 92606 297876 92612 297940
rect 92676 297938 92682 297940
rect 93577 297938 93643 297941
rect 92676 297936 93643 297938
rect 92676 297880 93582 297936
rect 93638 297880 93643 297936
rect 92676 297878 93643 297880
rect 92676 297876 92682 297878
rect 93577 297875 93643 297878
rect 94998 297876 95004 297940
rect 95068 297938 95074 297940
rect 95141 297938 95207 297941
rect 95068 297936 95207 297938
rect 95068 297880 95146 297936
rect 95202 297880 95207 297936
rect 95068 297878 95207 297880
rect 95558 297938 95618 298148
rect 95926 298074 95986 298148
rect 96521 298074 96587 298077
rect 96705 298076 96771 298077
rect 95926 298072 96587 298074
rect 95926 298016 96526 298072
rect 96582 298016 96587 298072
rect 95926 298014 96587 298016
rect 96521 298011 96587 298014
rect 96654 298012 96660 298076
rect 96724 298074 96771 298076
rect 97809 298074 97875 298077
rect 97942 298074 97948 298076
rect 96724 298072 96816 298074
rect 96766 298016 96816 298072
rect 96724 298014 96816 298016
rect 97809 298072 97948 298074
rect 97809 298016 97814 298072
rect 97870 298016 97948 298072
rect 97809 298014 97948 298016
rect 96724 298012 96771 298014
rect 96705 298011 96771 298012
rect 97809 298011 97875 298014
rect 97942 298012 97948 298014
rect 98012 298012 98018 298076
rect 99046 298012 99052 298076
rect 99116 298074 99122 298076
rect 99281 298074 99347 298077
rect 99116 298072 99347 298074
rect 99116 298016 99286 298072
rect 99342 298016 99347 298072
rect 99116 298014 99347 298016
rect 99116 298012 99122 298014
rect 99281 298011 99347 298014
rect 96429 297938 96495 297941
rect 95558 297936 96495 297938
rect 95558 297880 96434 297936
rect 96490 297880 96495 297936
rect 95558 297878 96495 297880
rect 95068 297876 95074 297878
rect 95141 297875 95207 297878
rect 96429 297875 96495 297878
rect 97022 297876 97028 297940
rect 97092 297938 97098 297940
rect 97717 297938 97783 297941
rect 97092 297936 97783 297938
rect 97092 297880 97722 297936
rect 97778 297880 97783 297936
rect 97092 297878 97783 297880
rect 97092 297876 97098 297878
rect 97717 297875 97783 297878
rect 98310 297876 98316 297940
rect 98380 297938 98386 297940
rect 99189 297938 99255 297941
rect 98380 297936 99255 297938
rect 98380 297880 99194 297936
rect 99250 297880 99255 297936
rect 98380 297878 99255 297880
rect 99422 297938 99482 298148
rect 100569 298076 100635 298077
rect 101857 298076 101923 298077
rect 100518 298074 100524 298076
rect 100478 298014 100524 298074
rect 100588 298072 100635 298076
rect 101806 298074 101812 298076
rect 100630 298016 100635 298072
rect 100518 298012 100524 298014
rect 100588 298012 100635 298016
rect 101766 298014 101812 298074
rect 101876 298072 101923 298076
rect 101918 298016 101923 298072
rect 101806 298012 101812 298014
rect 101876 298012 101923 298016
rect 102918 298074 102978 298148
rect 103237 298147 103303 298148
rect 103329 298074 103395 298077
rect 102918 298072 103395 298074
rect 102918 298016 103334 298072
rect 103390 298016 103395 298072
rect 102918 298014 103395 298016
rect 100569 298011 100635 298012
rect 101857 298011 101923 298012
rect 103329 298011 103395 298014
rect 104382 298012 104388 298076
rect 104452 298074 104458 298076
rect 104801 298074 104867 298077
rect 104452 298072 104867 298074
rect 104452 298016 104806 298072
rect 104862 298016 104867 298072
rect 104452 298014 104867 298016
rect 104452 298012 104458 298014
rect 104801 298011 104867 298014
rect 105670 298012 105676 298076
rect 105740 298074 105746 298076
rect 106181 298074 106247 298077
rect 105740 298072 106247 298074
rect 105740 298016 106186 298072
rect 106242 298016 106247 298072
rect 105740 298014 106247 298016
rect 105740 298012 105746 298014
rect 106181 298011 106247 298014
rect 106590 298012 106596 298076
rect 106660 298074 106666 298076
rect 106733 298074 106799 298077
rect 106660 298072 106799 298074
rect 106660 298016 106738 298072
rect 106794 298016 106799 298072
rect 106660 298014 106799 298016
rect 106660 298012 106666 298014
rect 106733 298011 106799 298014
rect 106958 298012 106964 298076
rect 107028 298074 107034 298076
rect 107469 298074 107535 298077
rect 107028 298072 107535 298074
rect 107028 298016 107474 298072
rect 107530 298016 107535 298072
rect 107028 298014 107535 298016
rect 107028 298012 107034 298014
rect 107469 298011 107535 298014
rect 107878 298012 107884 298076
rect 107948 298074 107954 298076
rect 108941 298074 109007 298077
rect 107948 298072 109007 298074
rect 107948 298016 108946 298072
rect 109002 298016 109007 298072
rect 107948 298014 109007 298016
rect 107948 298012 107954 298014
rect 108941 298011 109007 298014
rect 109350 298012 109356 298076
rect 109420 298074 109426 298076
rect 110321 298074 110387 298077
rect 109420 298072 110387 298074
rect 109420 298016 110326 298072
rect 110382 298016 110387 298072
rect 109420 298014 110387 298016
rect 109420 298012 109426 298014
rect 110321 298011 110387 298014
rect 110638 298012 110644 298076
rect 110708 298074 110714 298076
rect 111701 298074 111767 298077
rect 110708 298072 111767 298074
rect 110708 298016 111706 298072
rect 111762 298016 111767 298072
rect 110708 298014 111767 298016
rect 110708 298012 110714 298014
rect 111701 298011 111767 298014
rect 112989 298076 113055 298077
rect 112989 298072 113036 298076
rect 113100 298074 113106 298076
rect 112989 298016 112994 298072
rect 112989 298012 113036 298016
rect 113100 298014 113146 298074
rect 113100 298012 113106 298014
rect 114318 298012 114324 298076
rect 114388 298074 114394 298076
rect 114461 298074 114527 298077
rect 114388 298072 114527 298074
rect 114388 298016 114466 298072
rect 114522 298016 114527 298072
rect 114388 298014 114527 298016
rect 114388 298012 114394 298014
rect 112989 298011 113055 298012
rect 114461 298011 114527 298014
rect 115606 298012 115612 298076
rect 115676 298074 115682 298076
rect 115841 298074 115907 298077
rect 115676 298072 115907 298074
rect 115676 298016 115846 298072
rect 115902 298016 115907 298072
rect 115676 298014 115907 298016
rect 115676 298012 115682 298014
rect 115841 298011 115907 298014
rect 116894 298012 116900 298076
rect 116964 298074 116970 298076
rect 117221 298074 117287 298077
rect 116964 298072 117287 298074
rect 116964 298016 117226 298072
rect 117282 298016 117287 298072
rect 116964 298014 117287 298016
rect 116964 298012 116970 298014
rect 117221 298011 117287 298014
rect 215845 298076 215911 298077
rect 215845 298072 215892 298076
rect 215956 298074 215962 298076
rect 224953 298074 225019 298077
rect 225462 298074 225522 298148
rect 229142 298077 229202 298148
rect 258030 298077 258090 298150
rect 261518 298148 261524 298212
rect 261588 298148 261594 298212
rect 261886 298148 261892 298212
rect 261956 298148 261962 298212
rect 265198 298148 265204 298212
rect 265268 298148 265274 298212
rect 271822 298148 271828 298212
rect 271892 298148 271898 298212
rect 275502 298148 275508 298212
rect 275572 298148 275578 298212
rect 215845 298016 215850 298072
rect 215845 298012 215892 298016
rect 215956 298014 216002 298074
rect 224953 298072 225522 298074
rect 224953 298016 224958 298072
rect 225014 298016 225522 298072
rect 224953 298014 225522 298016
rect 226333 298074 226399 298077
rect 226742 298074 226748 298076
rect 226333 298072 226748 298074
rect 226333 298016 226338 298072
rect 226394 298016 226748 298072
rect 226333 298014 226748 298016
rect 215956 298012 215962 298014
rect 215845 298011 215911 298012
rect 224953 298011 225019 298014
rect 226333 298011 226399 298014
rect 226742 298012 226748 298014
rect 226812 298012 226818 298076
rect 227713 298074 227779 298077
rect 227846 298074 227852 298076
rect 227713 298072 227852 298074
rect 227713 298016 227718 298072
rect 227774 298016 227852 298072
rect 227713 298014 227852 298016
rect 227713 298011 227779 298014
rect 227846 298012 227852 298014
rect 227916 298012 227922 298076
rect 229142 298072 229251 298077
rect 229142 298016 229190 298072
rect 229246 298016 229251 298072
rect 229142 298014 229251 298016
rect 229185 298011 229251 298014
rect 230473 298074 230539 298077
rect 231342 298074 231348 298076
rect 230473 298072 231348 298074
rect 230473 298016 230478 298072
rect 230534 298016 231348 298072
rect 230473 298014 231348 298016
rect 230473 298011 230539 298014
rect 231342 298012 231348 298014
rect 231412 298012 231418 298076
rect 231853 298074 231919 298077
rect 232630 298074 232636 298076
rect 231853 298072 232636 298074
rect 231853 298016 231858 298072
rect 231914 298016 232636 298072
rect 231853 298014 232636 298016
rect 231853 298011 231919 298014
rect 232630 298012 232636 298014
rect 232700 298012 232706 298076
rect 233233 298074 233299 298077
rect 233550 298074 233556 298076
rect 233233 298072 233556 298074
rect 233233 298016 233238 298072
rect 233294 298016 233556 298072
rect 233233 298014 233556 298016
rect 233233 298011 233299 298014
rect 233550 298012 233556 298014
rect 233620 298012 233626 298076
rect 234613 298074 234679 298077
rect 237189 298076 237255 298077
rect 235022 298074 235028 298076
rect 234613 298072 235028 298074
rect 234613 298016 234618 298072
rect 234674 298016 235028 298072
rect 234613 298014 235028 298016
rect 234613 298011 234679 298014
rect 235022 298012 235028 298014
rect 235092 298012 235098 298076
rect 237189 298072 237236 298076
rect 237300 298074 237306 298076
rect 238753 298074 238819 298077
rect 239254 298074 239260 298076
rect 237189 298016 237194 298072
rect 237189 298012 237236 298016
rect 237300 298014 237346 298074
rect 238753 298072 239260 298074
rect 238753 298016 238758 298072
rect 238814 298016 239260 298072
rect 238753 298014 239260 298016
rect 237300 298012 237306 298014
rect 237189 298011 237255 298012
rect 238753 298011 238819 298014
rect 239254 298012 239260 298014
rect 239324 298012 239330 298076
rect 240133 298074 240199 298077
rect 240358 298074 240364 298076
rect 240133 298072 240364 298074
rect 240133 298016 240138 298072
rect 240194 298016 240364 298072
rect 240133 298014 240364 298016
rect 240133 298011 240199 298014
rect 240358 298012 240364 298014
rect 240428 298012 240434 298076
rect 240726 298012 240732 298076
rect 240796 298074 240802 298076
rect 241421 298074 241487 298077
rect 240796 298072 241487 298074
rect 240796 298016 241426 298072
rect 241482 298016 241487 298072
rect 240796 298014 241487 298016
rect 240796 298012 240802 298014
rect 241421 298011 241487 298014
rect 242893 298076 242959 298077
rect 244089 298076 244155 298077
rect 242893 298072 242940 298076
rect 243004 298074 243010 298076
rect 244038 298074 244044 298076
rect 242893 298016 242898 298072
rect 242893 298012 242940 298016
rect 243004 298014 243050 298074
rect 243998 298014 244044 298074
rect 244108 298072 244155 298076
rect 244150 298016 244155 298072
rect 243004 298012 243010 298014
rect 244038 298012 244044 298014
rect 244108 298012 244155 298016
rect 242893 298011 242959 298012
rect 244089 298011 244155 298012
rect 244273 298074 244339 298077
rect 245561 298076 245627 298077
rect 246849 298076 246915 298077
rect 244406 298074 244412 298076
rect 244273 298072 244412 298074
rect 244273 298016 244278 298072
rect 244334 298016 244412 298072
rect 244273 298014 244412 298016
rect 244273 298011 244339 298014
rect 244406 298012 244412 298014
rect 244476 298012 244482 298076
rect 245510 298074 245516 298076
rect 245470 298014 245516 298074
rect 245580 298072 245627 298076
rect 246798 298074 246804 298076
rect 245622 298016 245627 298072
rect 245510 298012 245516 298014
rect 245580 298012 245627 298016
rect 246758 298014 246804 298074
rect 246868 298072 246915 298076
rect 246910 298016 246915 298072
rect 246798 298012 246804 298014
rect 246868 298012 246915 298016
rect 247902 298012 247908 298076
rect 247972 298074 247978 298076
rect 248321 298074 248387 298077
rect 247972 298072 248387 298074
rect 247972 298016 248326 298072
rect 248382 298016 248387 298072
rect 247972 298014 248387 298016
rect 247972 298012 247978 298014
rect 245561 298011 245627 298012
rect 246849 298011 246915 298012
rect 248321 298011 248387 298014
rect 249374 298012 249380 298076
rect 249444 298074 249450 298076
rect 249701 298074 249767 298077
rect 249444 298072 249767 298074
rect 249444 298016 249706 298072
rect 249762 298016 249767 298072
rect 249444 298014 249767 298016
rect 249444 298012 249450 298014
rect 249701 298011 249767 298014
rect 250662 298012 250668 298076
rect 250732 298074 250738 298076
rect 251081 298074 251147 298077
rect 250732 298072 251147 298074
rect 250732 298016 251086 298072
rect 251142 298016 251147 298072
rect 250732 298014 251147 298016
rect 250732 298012 250738 298014
rect 251081 298011 251147 298014
rect 252369 298074 252435 298077
rect 252502 298074 252508 298076
rect 252369 298072 252508 298074
rect 252369 298016 252374 298072
rect 252430 298016 252508 298072
rect 252369 298014 252508 298016
rect 252369 298011 252435 298014
rect 252502 298012 252508 298014
rect 252572 298012 252578 298076
rect 253606 298012 253612 298076
rect 253676 298074 253682 298076
rect 253749 298074 253815 298077
rect 253676 298072 253815 298074
rect 253676 298016 253754 298072
rect 253810 298016 253815 298072
rect 253676 298014 253815 298016
rect 253676 298012 253682 298014
rect 253749 298011 253815 298014
rect 254894 298012 254900 298076
rect 254964 298074 254970 298076
rect 255129 298074 255195 298077
rect 254964 298072 255195 298074
rect 254964 298016 255134 298072
rect 255190 298016 255195 298072
rect 254964 298014 255195 298016
rect 254964 298012 254970 298014
rect 255129 298011 255195 298014
rect 255998 298012 256004 298076
rect 256068 298074 256074 298076
rect 256509 298074 256575 298077
rect 256068 298072 256575 298074
rect 256068 298016 256514 298072
rect 256570 298016 256575 298072
rect 256068 298014 256575 298016
rect 256068 298012 256074 298014
rect 256509 298011 256575 298014
rect 257102 298012 257108 298076
rect 257172 298074 257178 298076
rect 257797 298074 257863 298077
rect 257172 298072 257863 298074
rect 257172 298016 257802 298072
rect 257858 298016 257863 298072
rect 257172 298014 257863 298016
rect 257172 298012 257178 298014
rect 257797 298011 257863 298014
rect 257981 298072 258090 298077
rect 257981 298016 257986 298072
rect 258042 298016 258090 298072
rect 257981 298014 258090 298016
rect 259177 298074 259243 298077
rect 259310 298074 259316 298076
rect 259177 298072 259316 298074
rect 259177 298016 259182 298072
rect 259238 298016 259316 298072
rect 259177 298014 259316 298016
rect 257981 298011 258047 298014
rect 259177 298011 259243 298014
rect 259310 298012 259316 298014
rect 259380 298012 259386 298076
rect 260649 298074 260715 298077
rect 260782 298074 260788 298076
rect 260649 298072 260788 298074
rect 260649 298016 260654 298072
rect 260710 298016 260788 298072
rect 260649 298014 260788 298016
rect 260649 298011 260715 298014
rect 260782 298012 260788 298014
rect 260852 298012 260858 298076
rect 100661 297938 100727 297941
rect 99422 297936 100727 297938
rect 99422 297880 100666 297936
rect 100722 297880 100727 297936
rect 99422 297878 100727 297880
rect 98380 297876 98386 297878
rect 99189 297875 99255 297878
rect 100661 297875 100727 297878
rect 101438 297876 101444 297940
rect 101508 297938 101514 297940
rect 102041 297938 102107 297941
rect 101508 297936 102107 297938
rect 101508 297880 102046 297936
rect 102102 297880 102107 297936
rect 101508 297878 102107 297880
rect 101508 297876 101514 297878
rect 102041 297875 102107 297878
rect 104014 297876 104020 297940
rect 104084 297938 104090 297940
rect 104709 297938 104775 297941
rect 104084 297936 104775 297938
rect 104084 297880 104714 297936
rect 104770 297880 104775 297936
rect 104084 297878 104775 297880
rect 104084 297876 104090 297878
rect 104709 297875 104775 297878
rect 105302 297876 105308 297940
rect 105372 297938 105378 297940
rect 106089 297938 106155 297941
rect 105372 297936 106155 297938
rect 105372 297880 106094 297936
rect 106150 297880 106155 297936
rect 105372 297878 106155 297880
rect 105372 297876 105378 297878
rect 106089 297875 106155 297878
rect 107694 297876 107700 297940
rect 107764 297938 107770 297940
rect 108849 297938 108915 297941
rect 107764 297936 108915 297938
rect 107764 297880 108854 297936
rect 108910 297880 108915 297936
rect 107764 297878 108915 297880
rect 107764 297876 107770 297878
rect 108849 297875 108915 297878
rect 111926 297876 111932 297940
rect 111996 297938 112002 297940
rect 113081 297938 113147 297941
rect 111996 297936 113147 297938
rect 111996 297880 113086 297936
rect 113142 297880 113147 297936
rect 111996 297878 113147 297880
rect 111996 297876 112002 297878
rect 113081 297875 113147 297878
rect 237373 297938 237439 297941
rect 237782 297938 237788 297940
rect 237373 297936 237788 297938
rect 237373 297880 237378 297936
rect 237434 297880 237788 297936
rect 237373 297878 237788 297880
rect 237373 297875 237439 297878
rect 237782 297876 237788 297878
rect 237852 297876 237858 297940
rect 241513 297938 241579 297941
rect 242014 297938 242020 297940
rect 241513 297936 242020 297938
rect 241513 297880 241518 297936
rect 241574 297880 242020 297936
rect 241513 297878 242020 297880
rect 241513 297875 241579 297878
rect 242014 297876 242020 297878
rect 242084 297876 242090 297940
rect 243077 297938 243143 297941
rect 244181 297938 244247 297941
rect 243077 297936 244247 297938
rect 243077 297880 243082 297936
rect 243138 297880 244186 297936
rect 244242 297880 244247 297936
rect 243077 297878 244247 297880
rect 243077 297875 243143 297878
rect 244181 297875 244247 297878
rect 246614 297876 246620 297940
rect 246684 297938 246690 297940
rect 246757 297938 246823 297941
rect 246684 297936 246823 297938
rect 246684 297880 246762 297936
rect 246818 297880 246823 297936
rect 246684 297878 246823 297880
rect 246684 297876 246690 297878
rect 246757 297875 246823 297878
rect 247718 297876 247724 297940
rect 247788 297938 247794 297940
rect 248229 297938 248295 297941
rect 247788 297936 248295 297938
rect 247788 297880 248234 297936
rect 248290 297880 248295 297936
rect 247788 297878 248295 297880
rect 247788 297876 247794 297878
rect 248229 297875 248295 297878
rect 249006 297876 249012 297940
rect 249076 297938 249082 297940
rect 249609 297938 249675 297941
rect 249076 297936 249675 297938
rect 249076 297880 249614 297936
rect 249670 297880 249675 297936
rect 249076 297878 249675 297880
rect 249076 297876 249082 297878
rect 249609 297875 249675 297878
rect 250294 297876 250300 297940
rect 250364 297938 250370 297940
rect 250989 297938 251055 297941
rect 250364 297936 251055 297938
rect 250364 297880 250994 297936
rect 251050 297880 251055 297936
rect 250364 297878 251055 297880
rect 250364 297876 250370 297878
rect 250989 297875 251055 297878
rect 251398 297876 251404 297940
rect 251468 297938 251474 297940
rect 252277 297938 252343 297941
rect 251468 297936 252343 297938
rect 251468 297880 252282 297936
rect 252338 297880 252343 297936
rect 251468 297878 252343 297880
rect 251468 297876 251474 297878
rect 252277 297875 252343 297878
rect 253054 297876 253060 297940
rect 253124 297938 253130 297940
rect 253841 297938 253907 297941
rect 253124 297936 253907 297938
rect 253124 297880 253846 297936
rect 253902 297880 253907 297936
rect 253124 297878 253907 297880
rect 253124 297876 253130 297878
rect 253841 297875 253907 297878
rect 254526 297876 254532 297940
rect 254596 297938 254602 297940
rect 255221 297938 255287 297941
rect 254596 297936 255287 297938
rect 254596 297880 255226 297936
rect 255282 297880 255287 297936
rect 254596 297878 255287 297880
rect 254596 297876 254602 297878
rect 255221 297875 255287 297878
rect 255630 297876 255636 297940
rect 255700 297938 255706 297940
rect 256601 297938 256667 297941
rect 255700 297936 256667 297938
rect 255700 297880 256606 297936
rect 256662 297880 256667 297936
rect 255700 297878 256667 297880
rect 255700 297876 255706 297878
rect 256601 297875 256667 297878
rect 256734 297876 256740 297940
rect 256804 297938 256810 297940
rect 257889 297938 257955 297941
rect 256804 297936 257955 297938
rect 256804 297880 257894 297936
rect 257950 297880 257955 297936
rect 256804 297878 257955 297880
rect 256804 297876 256810 297878
rect 257889 297875 257955 297878
rect 259126 297876 259132 297940
rect 259196 297938 259202 297940
rect 259361 297938 259427 297941
rect 259196 297936 259427 297938
rect 259196 297880 259366 297936
rect 259422 297880 259427 297936
rect 259196 297878 259427 297880
rect 259196 297876 259202 297878
rect 259361 297875 259427 297878
rect 260598 297876 260604 297940
rect 260668 297938 260674 297940
rect 260741 297938 260807 297941
rect 260668 297936 260807 297938
rect 260668 297880 260746 297936
rect 260802 297880 260807 297936
rect 260668 297878 260807 297880
rect 261526 297938 261586 298148
rect 261894 298074 261954 298148
rect 262029 298074 262095 298077
rect 261894 298072 262095 298074
rect 261894 298016 262034 298072
rect 262090 298016 262095 298072
rect 261894 298014 262095 298016
rect 262029 298011 262095 298014
rect 263174 298012 263180 298076
rect 263244 298074 263250 298076
rect 263501 298074 263567 298077
rect 263244 298072 263567 298074
rect 263244 298016 263506 298072
rect 263562 298016 263567 298072
rect 263244 298014 263567 298016
rect 265206 298074 265266 298148
rect 266169 298074 266235 298077
rect 265206 298072 266235 298074
rect 265206 298016 266174 298072
rect 266230 298016 266235 298072
rect 265206 298014 266235 298016
rect 271830 298074 271890 298148
rect 273161 298074 273227 298077
rect 271830 298072 273227 298074
rect 271830 298016 273166 298072
rect 273222 298016 273227 298072
rect 271830 298014 273227 298016
rect 263244 298012 263250 298014
rect 263501 298011 263567 298014
rect 266169 298011 266235 298014
rect 273161 298011 273227 298014
rect 274398 298012 274404 298076
rect 274468 298074 274474 298076
rect 274541 298074 274607 298077
rect 274468 298072 274607 298074
rect 274468 298016 274546 298072
rect 274602 298016 274607 298072
rect 274468 298014 274607 298016
rect 275510 298074 275570 298148
rect 275921 298074 275987 298077
rect 275510 298072 275987 298074
rect 275510 298016 275926 298072
rect 275982 298016 275987 298072
rect 275510 298014 275987 298016
rect 274468 298012 274474 298014
rect 274541 298011 274607 298014
rect 275921 298011 275987 298014
rect 276790 298012 276796 298076
rect 276860 298074 276866 298076
rect 277301 298074 277367 298077
rect 276860 298072 277367 298074
rect 276860 298016 277306 298072
rect 277362 298016 277367 298072
rect 276860 298014 277367 298016
rect 276860 298012 276866 298014
rect 277301 298011 277367 298014
rect 262121 297938 262187 297941
rect 261526 297936 262187 297938
rect 261526 297880 262126 297936
rect 262182 297880 262187 297936
rect 261526 297878 262187 297880
rect 260668 297876 260674 297878
rect 260741 297875 260807 297878
rect 262121 297875 262187 297878
rect 262990 297876 262996 297940
rect 263060 297938 263066 297940
rect 263409 297938 263475 297941
rect 263060 297936 263475 297938
rect 263060 297880 263414 297936
rect 263470 297880 263475 297936
rect 263060 297878 263475 297880
rect 263060 297876 263066 297878
rect 263409 297875 263475 297878
rect 85798 297740 85804 297804
rect 85868 297802 85874 297804
rect 86861 297802 86927 297805
rect 85868 297800 86927 297802
rect 85868 297744 86866 297800
rect 86922 297744 86927 297800
rect 85868 297742 86927 297744
rect 85868 297740 85874 297742
rect 86861 297739 86927 297742
rect 100702 297740 100708 297804
rect 100772 297802 100778 297804
rect 101949 297802 102015 297805
rect 100772 297800 102015 297802
rect 100772 297744 101954 297800
rect 102010 297744 102015 297800
rect 100772 297742 102015 297744
rect 100772 297740 100778 297742
rect 101949 297739 102015 297742
rect 236494 297740 236500 297804
rect 236564 297802 236570 297804
rect 237281 297802 237347 297805
rect 236564 297800 237347 297802
rect 236564 297744 237286 297800
rect 237342 297744 237347 297800
rect 236564 297742 237347 297744
rect 236564 297740 236570 297742
rect 237281 297739 237347 297742
rect 241830 297740 241836 297804
rect 241900 297802 241906 297804
rect 242801 297802 242867 297805
rect 241900 297800 242867 297802
rect 241900 297744 242806 297800
rect 242862 297744 242867 297800
rect 241900 297742 242867 297744
rect 241900 297740 241906 297742
rect 242801 297739 242867 297742
rect 245694 297740 245700 297804
rect 245764 297802 245770 297804
rect 246941 297802 247007 297805
rect 245764 297800 247007 297802
rect 245764 297744 246946 297800
rect 247002 297744 247007 297800
rect 245764 297742 247007 297744
rect 245764 297740 245770 297742
rect 246941 297739 247007 297742
rect 251950 297740 251956 297804
rect 252020 297802 252026 297804
rect 252461 297802 252527 297805
rect 252020 297800 252527 297802
rect 252020 297744 252466 297800
rect 252522 297744 252527 297800
rect 252020 297742 252527 297744
rect 252020 297740 252026 297742
rect 252461 297739 252527 297742
rect 258390 297740 258396 297804
rect 258460 297802 258466 297804
rect 259269 297802 259335 297805
rect 258460 297800 259335 297802
rect 258460 297744 259274 297800
rect 259330 297744 259335 297800
rect 258460 297742 259335 297744
rect 258460 297740 258466 297742
rect 259269 297739 259335 297742
rect 267958 297468 267964 297532
rect 268028 297530 268034 297532
rect 269021 297530 269087 297533
rect 268028 297528 269087 297530
rect 268028 297472 269026 297528
rect 269082 297472 269087 297528
rect 268028 297470 269087 297472
rect 268028 297468 268034 297470
rect 269021 297467 269087 297470
rect 229461 297258 229527 297261
rect 230054 297258 230060 297260
rect 229461 297256 230060 297258
rect 229461 297200 229466 297256
rect 229522 297200 230060 297256
rect 229461 297198 230060 297200
rect 229461 297195 229527 297198
rect 230054 297196 230060 297198
rect 230124 297196 230130 297260
rect 83958 297060 83964 297124
rect 84028 297122 84034 297124
rect 85481 297122 85547 297125
rect 84028 297120 85547 297122
rect 84028 297064 85486 297120
rect 85542 297064 85547 297120
rect 84028 297062 85547 297064
rect 84028 297060 84034 297062
rect 85481 297059 85547 297062
rect 238661 297122 238727 297125
rect 240041 297122 240107 297125
rect 238661 297120 240107 297122
rect 238661 297064 238666 297120
rect 238722 297064 240046 297120
rect 240102 297064 240107 297120
rect 238661 297062 240107 297064
rect 238661 297059 238727 297062
rect 240041 297059 240107 297062
rect 266670 297060 266676 297124
rect 266740 297122 266746 297124
rect 267549 297122 267615 297125
rect 266740 297120 267615 297122
rect 266740 297064 267554 297120
rect 267610 297064 267615 297120
rect 266740 297062 267615 297064
rect 266740 297060 266746 297062
rect 267549 297059 267615 297062
rect 264094 296924 264100 296988
rect 264164 296986 264170 296988
rect 264789 296986 264855 296989
rect 264164 296984 264855 296986
rect 264164 296928 264794 296984
rect 264850 296928 264855 296984
rect 264164 296926 264855 296928
rect 264164 296924 264170 296926
rect 264789 296923 264855 296926
rect 266854 296924 266860 296988
rect 266924 296986 266930 296988
rect 267641 296986 267707 296989
rect 266924 296984 267707 296986
rect 266924 296928 267646 296984
rect 267702 296928 267707 296984
rect 266924 296926 267707 296928
rect 266924 296924 266930 296926
rect 267641 296923 267707 296926
rect 238334 296788 238340 296852
rect 238404 296850 238410 296852
rect 238661 296850 238727 296853
rect 238404 296848 238727 296850
rect 238404 296792 238666 296848
rect 238722 296792 238727 296848
rect 238404 296790 238727 296792
rect 238404 296788 238410 296790
rect 238661 296787 238727 296790
rect 264462 296788 264468 296852
rect 264532 296850 264538 296852
rect 264881 296850 264947 296853
rect 264532 296848 264947 296850
rect 264532 296792 264886 296848
rect 264942 296792 264947 296848
rect 264532 296790 264947 296792
rect 264532 296788 264538 296790
rect 264881 296787 264947 296790
rect 265750 296788 265756 296852
rect 265820 296850 265826 296852
rect 266261 296850 266327 296853
rect 265820 296848 266327 296850
rect 265820 296792 266266 296848
rect 266322 296792 266327 296848
rect 265820 296790 266327 296792
rect 265820 296788 265826 296790
rect 266261 296787 266327 296790
rect 267457 296850 267523 296853
rect 267590 296850 267596 296852
rect 267457 296848 267596 296850
rect 267457 296792 267462 296848
rect 267518 296792 267596 296848
rect 267457 296790 267596 296792
rect 267457 296787 267523 296790
rect 267590 296788 267596 296790
rect 267660 296788 267666 296852
rect 269246 296788 269252 296852
rect 269316 296850 269322 296852
rect 270401 296850 270467 296853
rect 269316 296848 270467 296850
rect 269316 296792 270406 296848
rect 270462 296792 270467 296848
rect 269316 296790 270467 296792
rect 269316 296788 269322 296790
rect 270401 296787 270467 296790
rect 270534 296788 270540 296852
rect 270604 296850 270610 296852
rect 271781 296850 271847 296853
rect 270604 296848 271847 296850
rect 270604 296792 271786 296848
rect 271842 296792 271847 296848
rect 270604 296790 271847 296792
rect 270604 296788 270610 296790
rect 271781 296787 271847 296790
rect 273069 296852 273135 296853
rect 273069 296848 273116 296852
rect 273180 296850 273186 296852
rect 273069 296792 273074 296848
rect 273069 296788 273116 296792
rect 273180 296790 273226 296850
rect 273180 296788 273186 296790
rect 273069 296787 273135 296788
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 408493 249658 408559 249661
rect 408493 249656 409338 249658
rect 408493 249600 408498 249656
rect 408554 249600 409338 249656
rect 408493 249598 409338 249600
rect 408493 249595 408559 249598
rect 187601 249522 187667 249525
rect 187601 249520 190164 249522
rect 187601 249464 187606 249520
rect 187662 249464 190164 249520
rect 187601 249462 190164 249464
rect 187601 249459 187667 249462
rect 409278 249084 409338 249598
rect 187509 248434 187575 248437
rect 187509 248432 189826 248434
rect 187509 248376 187514 248432
rect 187570 248406 189826 248432
rect 187570 248376 190010 248406
rect 187509 248374 190010 248376
rect 187509 248371 187575 248374
rect 189766 248366 190010 248374
rect 189766 248346 190072 248366
rect 189950 248306 190072 248346
rect 409321 247754 409387 247757
rect 409321 247752 409522 247754
rect 409321 247696 409326 247752
rect 409382 247696 409522 247752
rect 409321 247694 409522 247696
rect 409321 247691 409387 247694
rect 187601 247346 187667 247349
rect 187601 247344 189642 247346
rect 187601 247288 187606 247344
rect 187662 247318 189642 247344
rect 187662 247288 190164 247318
rect 187601 247286 190164 247288
rect 187601 247283 187667 247286
rect 189582 247258 190164 247286
rect 409462 247180 409522 247694
rect 187325 246122 187391 246125
rect 187325 246120 189642 246122
rect 187325 246064 187330 246120
rect 187386 246094 189642 246120
rect 187386 246064 190164 246094
rect 187325 246062 190164 246064
rect 187325 246059 187391 246062
rect 189582 246034 190164 246062
rect 583520 245428 584960 245668
rect 411253 245170 411319 245173
rect 409860 245168 411319 245170
rect 409860 245112 411258 245168
rect 411314 245112 411319 245168
rect 409860 245110 411319 245112
rect 411253 245107 411319 245110
rect 187601 245034 187667 245037
rect 187601 245032 189642 245034
rect 187601 244976 187606 245032
rect 187662 245006 189642 245032
rect 187662 244976 190164 245006
rect 187601 244974 190164 244976
rect 187601 244971 187667 244974
rect 189582 244946 190164 244974
rect 186313 243946 186379 243949
rect 186313 243944 189642 243946
rect 186313 243888 186318 243944
rect 186374 243918 189642 243944
rect 186374 243888 190164 243918
rect 186313 243886 190164 243888
rect 186313 243883 186379 243886
rect 189582 243858 190164 243886
rect 410517 243266 410583 243269
rect 409860 243264 410583 243266
rect 409860 243208 410522 243264
rect 410578 243208 410583 243264
rect 409860 243206 410583 243208
rect 410517 243203 410583 243206
rect 186313 242722 186379 242725
rect 186313 242720 189642 242722
rect 186313 242664 186318 242720
rect 186374 242694 189642 242720
rect 186374 242664 190164 242694
rect 186313 242662 190164 242664
rect 186313 242659 186379 242662
rect 189582 242634 190164 242662
rect 186405 241634 186471 241637
rect 186405 241632 189642 241634
rect 186405 241576 186410 241632
rect 186466 241606 189642 241632
rect 186466 241576 190164 241606
rect 186405 241574 190164 241576
rect 186405 241571 186471 241574
rect 189582 241546 190164 241574
rect 410425 241226 410491 241229
rect 409860 241224 410491 241226
rect -960 240940 480 241180
rect 409860 241168 410430 241224
rect 410486 241168 410491 241224
rect 409860 241166 410491 241168
rect 410425 241163 410491 241166
rect 186313 240546 186379 240549
rect 186313 240544 189642 240546
rect 186313 240488 186318 240544
rect 186374 240518 189642 240544
rect 186374 240488 190164 240518
rect 186313 240486 190164 240488
rect 186313 240483 186379 240486
rect 189582 240458 190164 240486
rect 186313 239458 186379 239461
rect 186313 239456 189642 239458
rect 186313 239400 186318 239456
rect 186374 239430 189642 239456
rect 186374 239400 190164 239430
rect 186313 239398 190164 239400
rect 186313 239395 186379 239398
rect 189582 239370 190164 239398
rect 411621 239322 411687 239325
rect 409860 239320 411687 239322
rect 409860 239264 411626 239320
rect 411682 239264 411687 239320
rect 409860 239262 411687 239264
rect 411621 239259 411687 239262
rect 186313 238234 186379 238237
rect 186313 238232 189642 238234
rect 186313 238176 186318 238232
rect 186374 238206 189642 238232
rect 186374 238176 190164 238206
rect 186313 238174 190164 238176
rect 186313 238171 186379 238174
rect 189582 238146 190164 238174
rect 411529 237282 411595 237285
rect 409860 237280 411595 237282
rect 409860 237224 411534 237280
rect 411590 237224 411595 237280
rect 409860 237222 411595 237224
rect 411529 237219 411595 237222
rect 186313 237146 186379 237149
rect 186313 237144 189642 237146
rect 186313 237088 186318 237144
rect 186374 237118 189642 237144
rect 186374 237088 190164 237118
rect 186313 237086 190164 237088
rect 186313 237083 186379 237086
rect 189582 237058 190164 237086
rect 186405 236058 186471 236061
rect 186405 236056 189642 236058
rect 186405 236000 186410 236056
rect 186466 236030 189642 236056
rect 186466 236000 190164 236030
rect 186405 235998 190164 236000
rect 186405 235995 186471 235998
rect 189582 235970 190164 235998
rect 411253 235378 411319 235381
rect 409860 235376 411319 235378
rect 409860 235320 411258 235376
rect 411314 235320 411319 235376
rect 409860 235318 411319 235320
rect 411253 235315 411319 235318
rect 186313 234834 186379 234837
rect 186313 234832 189642 234834
rect 186313 234776 186318 234832
rect 186374 234806 189642 234832
rect 186374 234776 190164 234806
rect 186313 234774 190164 234776
rect 186313 234771 186379 234774
rect 189582 234746 190164 234774
rect 186313 233746 186379 233749
rect 409321 233746 409387 233749
rect 186313 233744 189642 233746
rect 186313 233688 186318 233744
rect 186374 233718 189642 233744
rect 409278 233744 409387 233746
rect 186374 233688 190164 233718
rect 186313 233686 190164 233688
rect 186313 233683 186379 233686
rect 189582 233658 190164 233686
rect 409278 233688 409326 233744
rect 409382 233688 409387 233744
rect 409278 233683 409387 233688
rect 409278 233308 409338 233683
rect 186313 232658 186379 232661
rect 186313 232656 189642 232658
rect 186313 232600 186318 232656
rect 186374 232630 189642 232656
rect 186374 232600 190164 232630
rect 186313 232598 190164 232600
rect 186313 232595 186379 232598
rect 189582 232570 190164 232598
rect 579613 232386 579679 232389
rect 583520 232386 584960 232476
rect 579613 232384 584960 232386
rect 579613 232328 579618 232384
rect 579674 232328 584960 232384
rect 579613 232326 584960 232328
rect 579613 232323 579679 232326
rect 583520 232236 584960 232326
rect 409321 231842 409387 231845
rect 409321 231840 409522 231842
rect 409321 231784 409326 231840
rect 409382 231784 409522 231840
rect 409321 231782 409522 231784
rect 409321 231779 409387 231782
rect 186313 231434 186379 231437
rect 186313 231432 189642 231434
rect 186313 231376 186318 231432
rect 186374 231406 189642 231432
rect 186374 231376 190164 231406
rect 409462 231404 409522 231782
rect 186313 231374 190164 231376
rect 186313 231371 186379 231374
rect 189582 231346 190164 231374
rect 409321 230074 409387 230077
rect 409278 230072 409387 230074
rect 409278 230016 409326 230072
rect 409382 230016 409387 230072
rect 409278 230011 409387 230016
rect 409278 229500 409338 230011
rect 186313 229258 186379 229261
rect 186313 229256 189642 229258
rect 186313 229200 186318 229256
rect 186374 229230 189642 229256
rect 186374 229200 190164 229230
rect 186313 229198 190164 229200
rect 186313 229195 186379 229198
rect 189582 229170 190164 229198
rect 186313 228170 186379 228173
rect 186313 228168 189642 228170
rect -960 227884 480 228124
rect 186313 228112 186318 228168
rect 186374 228142 189642 228168
rect 186374 228112 190164 228142
rect 186313 228110 190164 228112
rect 186313 228107 186379 228110
rect 189582 228082 190164 228110
rect 410333 227490 410399 227493
rect 409860 227488 410399 227490
rect 409860 227432 410338 227488
rect 410394 227432 410399 227488
rect 409860 227430 410399 227432
rect 410333 227427 410399 227430
rect 410057 226130 410123 226133
rect 409830 226128 410123 226130
rect 409830 226072 410062 226128
rect 410118 226072 410123 226128
rect 409830 226070 410123 226072
rect 189398 225730 190072 225790
rect 186681 225722 186747 225725
rect 189398 225722 189458 225730
rect 186681 225720 189458 225722
rect 186681 225664 186686 225720
rect 186742 225664 189458 225720
rect 186681 225662 189458 225664
rect 186681 225659 186747 225662
rect 409830 225556 409890 226070
rect 410057 226067 410123 226070
rect 187509 224770 187575 224773
rect 187509 224768 189642 224770
rect 187509 224712 187514 224768
rect 187570 224742 189642 224768
rect 187570 224712 190164 224742
rect 187509 224710 190164 224712
rect 187509 224707 187575 224710
rect 189582 224682 190164 224710
rect 187601 223546 187667 223549
rect 187601 223544 189642 223546
rect 187601 223488 187606 223544
rect 187662 223518 189642 223544
rect 187662 223488 190164 223518
rect 187601 223486 190164 223488
rect 187601 223483 187667 223486
rect 189582 223458 190164 223486
rect 409830 223274 409890 223516
rect 409965 223274 410031 223277
rect 409830 223272 410031 223274
rect 409830 223216 409970 223272
rect 410026 223216 410031 223272
rect 409830 223214 410031 223216
rect 409965 223211 410031 223214
rect 189398 222330 190072 222390
rect 186313 222322 186379 222325
rect 189398 222322 189458 222330
rect 186313 222320 189458 222322
rect 186313 222264 186318 222320
rect 186374 222264 189458 222320
rect 186313 222262 189458 222264
rect 186313 222259 186379 222262
rect 410241 221642 410307 221645
rect 409860 221640 410307 221642
rect 409860 221584 410246 221640
rect 410302 221584 410307 221640
rect 409860 221582 410307 221584
rect 410241 221579 410307 221582
rect 189398 221242 190072 221302
rect 186313 221234 186379 221237
rect 189398 221234 189458 221242
rect 186313 221232 189458 221234
rect 186313 221176 186318 221232
rect 186374 221176 189458 221232
rect 186313 221174 189458 221176
rect 186313 221171 186379 221174
rect 189398 220018 190072 220078
rect 186313 220010 186379 220013
rect 189398 220010 189458 220018
rect 186313 220008 189458 220010
rect 186313 219952 186318 220008
rect 186374 219952 189458 220008
rect 186313 219950 189458 219952
rect 186313 219947 186379 219950
rect 411713 219602 411779 219605
rect 409860 219600 411779 219602
rect 409860 219544 411718 219600
rect 411774 219544 411779 219600
rect 409860 219542 411779 219544
rect 411713 219539 411779 219542
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 189398 218930 190072 218990
rect 186313 218922 186379 218925
rect 189398 218922 189458 218930
rect 186313 218920 189458 218922
rect 186313 218864 186318 218920
rect 186374 218864 189458 218920
rect 583520 218908 584960 218998
rect 186313 218862 189458 218864
rect 186313 218859 186379 218862
rect 189398 217842 190072 217902
rect 186405 217834 186471 217837
rect 189398 217834 189458 217842
rect 186405 217832 189458 217834
rect 186405 217776 186410 217832
rect 186466 217776 189458 217832
rect 186405 217774 189458 217776
rect 186405 217771 186471 217774
rect 410149 217698 410215 217701
rect 409860 217696 410215 217698
rect 409860 217640 410154 217696
rect 410210 217640 410215 217696
rect 409860 217638 410215 217640
rect 410149 217635 410215 217638
rect 189398 216754 190072 216814
rect 186313 216746 186379 216749
rect 189398 216746 189458 216754
rect 186313 216744 189458 216746
rect 186313 216688 186318 216744
rect 186374 216688 189458 216744
rect 186313 216686 189458 216688
rect 186313 216683 186379 216686
rect 411437 215658 411503 215661
rect 409860 215656 411503 215658
rect 409860 215600 411442 215656
rect 411498 215600 411503 215656
rect 409860 215598 411503 215600
rect 411437 215595 411503 215598
rect 189398 215530 190072 215590
rect 186313 215522 186379 215525
rect 189398 215522 189458 215530
rect 186313 215520 189458 215522
rect 186313 215464 186318 215520
rect 186374 215464 189458 215520
rect 186313 215462 189458 215464
rect 186313 215459 186379 215462
rect -960 214828 480 215068
rect 189398 214442 190072 214502
rect 186313 214434 186379 214437
rect 189398 214434 189458 214442
rect 186313 214432 189458 214434
rect 186313 214376 186318 214432
rect 186374 214376 189458 214432
rect 186313 214374 189458 214376
rect 186313 214371 186379 214374
rect 411345 213754 411411 213757
rect 409860 213752 411411 213754
rect 409860 213696 411350 213752
rect 411406 213696 411411 213752
rect 409860 213694 411411 213696
rect 411345 213691 411411 213694
rect 189398 213354 190072 213414
rect 186313 213346 186379 213349
rect 189398 213346 189458 213354
rect 186313 213344 189458 213346
rect 186313 213288 186318 213344
rect 186374 213288 189458 213344
rect 186313 213286 189458 213288
rect 186313 213283 186379 213286
rect 409873 212394 409939 212397
rect 409830 212392 409939 212394
rect 409830 212336 409878 212392
rect 409934 212336 409939 212392
rect 409830 212331 409939 212336
rect 189398 212130 190072 212190
rect 186957 212122 187023 212125
rect 189398 212122 189458 212130
rect 186957 212120 189458 212122
rect 186957 212064 186962 212120
rect 187018 212064 189458 212120
rect 186957 212062 189458 212064
rect 186957 212059 187023 212062
rect 409830 211820 409890 212331
rect 186313 211170 186379 211173
rect 186313 211168 189826 211170
rect 186313 211112 186318 211168
rect 186374 211142 189826 211168
rect 186374 211112 190010 211142
rect 186313 211110 190010 211112
rect 186313 211107 186379 211110
rect 189766 211102 190010 211110
rect 189766 211082 190072 211102
rect 189950 211042 190072 211082
rect 189398 209954 190072 210014
rect 186313 209946 186379 209949
rect 189398 209946 189458 209954
rect 186313 209944 189458 209946
rect 186313 209888 186318 209944
rect 186374 209888 189458 209944
rect 186313 209886 189458 209888
rect 186313 209883 186379 209886
rect 411253 209810 411319 209813
rect 409860 209808 411319 209810
rect 409860 209752 411258 209808
rect 411314 209752 411319 209808
rect 409860 209750 411319 209752
rect 411253 209747 411319 209750
rect 189398 208730 190072 208790
rect 186313 208722 186379 208725
rect 189398 208722 189458 208730
rect 186313 208720 189458 208722
rect 186313 208664 186318 208720
rect 186374 208664 189458 208720
rect 186313 208662 189458 208664
rect 186313 208659 186379 208662
rect 411253 207906 411319 207909
rect 409860 207904 411319 207906
rect 409860 207848 411258 207904
rect 411314 207848 411319 207904
rect 409860 207846 411319 207848
rect 411253 207843 411319 207846
rect 189398 207642 190072 207702
rect 186313 207634 186379 207637
rect 189398 207634 189458 207642
rect 186313 207632 189458 207634
rect 186313 207576 186318 207632
rect 186374 207576 189458 207632
rect 186313 207574 189458 207576
rect 186313 207571 186379 207574
rect 189398 206554 190072 206614
rect 186313 206546 186379 206549
rect 189398 206546 189458 206554
rect 186313 206544 189458 206546
rect 186313 206488 186318 206544
rect 186374 206488 189458 206544
rect 186313 206486 189458 206488
rect 186313 206483 186379 206486
rect 411253 205866 411319 205869
rect 409860 205864 411319 205866
rect 409860 205808 411258 205864
rect 411314 205808 411319 205864
rect 409860 205806 411319 205808
rect 411253 205803 411319 205806
rect 583520 205580 584960 205820
rect 189398 205466 190072 205526
rect 187049 205458 187115 205461
rect 189398 205458 189458 205466
rect 187049 205456 189458 205458
rect 187049 205400 187054 205456
rect 187110 205400 189458 205456
rect 187049 205398 189458 205400
rect 187049 205395 187115 205398
rect 186313 204370 186379 204373
rect 186313 204368 189642 204370
rect 186313 204312 186318 204368
rect 186374 204342 189642 204368
rect 186374 204312 190164 204342
rect 186313 204310 190164 204312
rect 186313 204307 186379 204310
rect 189582 204282 190164 204310
rect 411253 203962 411319 203965
rect 409860 203960 411319 203962
rect 409860 203904 411258 203960
rect 411314 203904 411319 203960
rect 409860 203902 411319 203904
rect 411253 203899 411319 203902
rect 189398 203154 190072 203214
rect 186313 203146 186379 203149
rect 189398 203146 189458 203154
rect 186313 203144 189458 203146
rect 186313 203088 186318 203144
rect 186374 203088 189458 203144
rect 186313 203086 189458 203088
rect 186313 203083 186379 203086
rect 189398 202066 190072 202126
rect 186313 202058 186379 202061
rect 189398 202058 189458 202066
rect 186313 202056 189458 202058
rect -960 201772 480 202012
rect 186313 202000 186318 202056
rect 186374 202000 189458 202056
rect 186313 201998 189458 202000
rect 186313 201995 186379 201998
rect 411897 201922 411963 201925
rect 409860 201920 411963 201922
rect 409860 201864 411902 201920
rect 411958 201864 411963 201920
rect 409860 201862 411963 201864
rect 411897 201859 411963 201862
rect 189398 200842 190072 200902
rect 186313 200834 186379 200837
rect 189398 200834 189458 200842
rect 186313 200832 189458 200834
rect 186313 200776 186318 200832
rect 186374 200776 189458 200832
rect 186313 200774 189458 200776
rect 186313 200771 186379 200774
rect 412081 200018 412147 200021
rect 409860 200016 412147 200018
rect 409860 199960 412086 200016
rect 412142 199960 412147 200016
rect 409860 199958 412147 199960
rect 412081 199955 412147 199958
rect 189398 199754 190072 199814
rect 186405 199746 186471 199749
rect 189398 199746 189458 199754
rect 186405 199744 189458 199746
rect 186405 199688 186410 199744
rect 186466 199688 189458 199744
rect 186405 199686 189458 199688
rect 186405 199683 186471 199686
rect 186313 198794 186379 198797
rect 186313 198792 189642 198794
rect 186313 198736 186318 198792
rect 186374 198766 189642 198792
rect 186374 198736 190164 198766
rect 186313 198734 190164 198736
rect 186313 198731 186379 198734
rect 189582 198706 190164 198734
rect 411253 197978 411319 197981
rect 409860 197976 411319 197978
rect 409860 197920 411258 197976
rect 411314 197920 411319 197976
rect 409860 197918 411319 197920
rect 411253 197915 411319 197918
rect 189398 197578 190072 197638
rect 186313 197570 186379 197573
rect 189398 197570 189458 197578
rect 186313 197568 189458 197570
rect 186313 197512 186318 197568
rect 186374 197512 189458 197568
rect 186313 197510 189458 197512
rect 186313 197507 186379 197510
rect 189398 196354 190072 196414
rect 186313 196346 186379 196349
rect 189398 196346 189458 196354
rect 186313 196344 189458 196346
rect 186313 196288 186318 196344
rect 186374 196288 189458 196344
rect 186313 196286 189458 196288
rect 186313 196283 186379 196286
rect 411253 196074 411319 196077
rect 409860 196072 411319 196074
rect 409860 196016 411258 196072
rect 411314 196016 411319 196072
rect 409860 196014 411319 196016
rect 411253 196011 411319 196014
rect 189398 195266 190072 195326
rect 186313 195258 186379 195261
rect 189398 195258 189458 195266
rect 186313 195256 189458 195258
rect 186313 195200 186318 195256
rect 186374 195200 189458 195256
rect 186313 195198 189458 195200
rect 186313 195195 186379 195198
rect 189398 194178 190072 194238
rect 186313 194170 186379 194173
rect 189398 194170 189458 194178
rect 411989 194170 412055 194173
rect 186313 194168 189458 194170
rect 186313 194112 186318 194168
rect 186374 194112 189458 194168
rect 186313 194110 189458 194112
rect 409860 194168 412055 194170
rect 409860 194112 411994 194168
rect 412050 194112 412055 194168
rect 409860 194110 412055 194112
rect 186313 194107 186379 194110
rect 411989 194107 412055 194110
rect 189398 192954 190072 193014
rect 186405 192946 186471 192949
rect 189398 192946 189458 192954
rect 186405 192944 189458 192946
rect 186405 192888 186410 192944
rect 186466 192888 189458 192944
rect 186405 192886 189458 192888
rect 186405 192883 186471 192886
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 411253 192130 411319 192133
rect 409860 192128 411319 192130
rect 409860 192072 411258 192128
rect 411314 192072 411319 192128
rect 409860 192070 411319 192072
rect 411253 192067 411319 192070
rect 189398 191866 190072 191926
rect 186313 191858 186379 191861
rect 189398 191858 189458 191866
rect 186313 191856 189458 191858
rect 186313 191800 186318 191856
rect 186374 191800 189458 191856
rect 186313 191798 189458 191800
rect 186313 191795 186379 191798
rect 189398 190778 190072 190838
rect 186313 190770 186379 190773
rect 189398 190770 189458 190778
rect 186313 190768 189458 190770
rect 186313 190712 186318 190768
rect 186374 190712 189458 190768
rect 186313 190710 189458 190712
rect 186313 190707 186379 190710
rect 411253 190226 411319 190229
rect 409860 190224 411319 190226
rect 409860 190168 411258 190224
rect 411314 190168 411319 190224
rect 409860 190166 411319 190168
rect 411253 190163 411319 190166
rect 189398 189554 190072 189614
rect 186313 189546 186379 189549
rect 189398 189546 189458 189554
rect 186313 189544 189458 189546
rect 186313 189488 186318 189544
rect 186374 189488 189458 189544
rect 186313 189486 189458 189488
rect 186313 189483 186379 189486
rect -960 188716 480 188956
rect 189398 188466 190072 188526
rect 186313 188458 186379 188461
rect 189398 188458 189458 188466
rect 186313 188456 189458 188458
rect 186313 188400 186318 188456
rect 186374 188400 189458 188456
rect 186313 188398 189458 188400
rect 186313 188395 186379 188398
rect 411253 188186 411319 188189
rect 409860 188184 411319 188186
rect 409860 188128 411258 188184
rect 411314 188128 411319 188184
rect 409860 188126 411319 188128
rect 411253 188123 411319 188126
rect 189398 187378 190072 187438
rect 186405 187370 186471 187373
rect 189398 187370 189458 187378
rect 186405 187368 189458 187370
rect 186405 187312 186410 187368
rect 186466 187312 189458 187368
rect 186405 187310 189458 187312
rect 186405 187307 186471 187310
rect 186313 186418 186379 186421
rect 186313 186416 189642 186418
rect 186313 186360 186318 186416
rect 186374 186390 189642 186416
rect 186374 186360 190164 186390
rect 186313 186358 190164 186360
rect 186313 186355 186379 186358
rect 189582 186330 190164 186358
rect 411253 186282 411319 186285
rect 409860 186280 411319 186282
rect 409860 186224 411258 186280
rect 411314 186224 411319 186280
rect 409860 186222 411319 186224
rect 411253 186219 411319 186222
rect 189398 185066 190072 185126
rect 187141 185058 187207 185061
rect 189398 185058 189458 185066
rect 187141 185056 189458 185058
rect 187141 185000 187146 185056
rect 187202 185000 189458 185056
rect 187141 184998 189458 185000
rect 187141 184995 187207 184998
rect 411253 184242 411319 184245
rect 409860 184240 411319 184242
rect 409860 184184 411258 184240
rect 411314 184184 411319 184240
rect 409860 184182 411319 184184
rect 411253 184179 411319 184182
rect 189398 183978 190072 184038
rect 186313 183970 186379 183973
rect 189398 183970 189458 183978
rect 186313 183968 189458 183970
rect 186313 183912 186318 183968
rect 186374 183912 189458 183968
rect 186313 183910 189458 183912
rect 186313 183907 186379 183910
rect 189398 182890 190072 182950
rect 186313 182882 186379 182885
rect 189398 182882 189458 182890
rect 186313 182880 189458 182882
rect 186313 182824 186318 182880
rect 186374 182824 189458 182880
rect 186313 182822 189458 182824
rect 186313 182819 186379 182822
rect 411253 182338 411319 182341
rect 409860 182336 411319 182338
rect 409860 182280 411258 182336
rect 411314 182280 411319 182336
rect 409860 182278 411319 182280
rect 411253 182275 411319 182278
rect 189398 181666 190072 181726
rect 186313 181658 186379 181661
rect 189398 181658 189458 181666
rect 186313 181656 189458 181658
rect 186313 181600 186318 181656
rect 186374 181600 189458 181656
rect 186313 181598 189458 181600
rect 186313 181595 186379 181598
rect 189398 180578 190072 180638
rect 186405 180570 186471 180573
rect 189398 180570 189458 180578
rect 186405 180568 189458 180570
rect 186405 180512 186410 180568
rect 186466 180512 189458 180568
rect 186405 180510 189458 180512
rect 186405 180507 186471 180510
rect 411253 180298 411319 180301
rect 409860 180296 411319 180298
rect 409860 180240 411258 180296
rect 411314 180240 411319 180296
rect 409860 180238 411319 180240
rect 411253 180235 411319 180238
rect 189398 179490 190072 179550
rect 186313 179482 186379 179485
rect 189398 179482 189458 179490
rect 186313 179480 189458 179482
rect 186313 179424 186318 179480
rect 186374 179424 189458 179480
rect 186313 179422 189458 179424
rect 186313 179419 186379 179422
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 411253 178394 411319 178397
rect 409860 178392 411319 178394
rect 409860 178336 411258 178392
rect 411314 178336 411319 178392
rect 409860 178334 411319 178336
rect 411253 178331 411319 178334
rect 189398 178266 190072 178326
rect 186313 178258 186379 178261
rect 189398 178258 189458 178266
rect 186313 178256 189458 178258
rect 186313 178200 186318 178256
rect 186374 178200 189458 178256
rect 186313 178198 189458 178200
rect 186313 178195 186379 178198
rect 189398 177178 190072 177238
rect 186313 177170 186379 177173
rect 189398 177170 189458 177178
rect 186313 177168 189458 177170
rect 186313 177112 186318 177168
rect 186374 177112 189458 177168
rect 186313 177110 189458 177112
rect 186313 177107 186379 177110
rect 411253 176490 411319 176493
rect 409860 176488 411319 176490
rect 409860 176432 411258 176488
rect 411314 176432 411319 176488
rect 409860 176430 411319 176432
rect 411253 176427 411319 176430
rect 189398 176090 190072 176150
rect 186313 176082 186379 176085
rect 189398 176082 189458 176090
rect 186313 176080 189458 176082
rect -960 175796 480 176036
rect 186313 176024 186318 176080
rect 186374 176024 189458 176080
rect 186313 176022 189458 176024
rect 186313 176019 186379 176022
rect 189398 175002 190072 175062
rect 186313 174994 186379 174997
rect 189398 174994 189458 175002
rect 186313 174992 189458 174994
rect 186313 174936 186318 174992
rect 186374 174936 189458 174992
rect 186313 174934 189458 174936
rect 186313 174931 186379 174934
rect 411253 174450 411319 174453
rect 409860 174448 411319 174450
rect 409860 174392 411258 174448
rect 411314 174392 411319 174448
rect 409860 174390 411319 174392
rect 411253 174387 411319 174390
rect 189398 173778 190072 173838
rect 187233 173770 187299 173773
rect 189398 173770 189458 173778
rect 187233 173768 189458 173770
rect 187233 173712 187238 173768
rect 187294 173712 189458 173768
rect 187233 173710 189458 173712
rect 187233 173707 187299 173710
rect 189398 172690 190072 172750
rect 186313 172682 186379 172685
rect 189398 172682 189458 172690
rect 186313 172680 189458 172682
rect 186313 172624 186318 172680
rect 186374 172624 189458 172680
rect 186313 172622 189458 172624
rect 186313 172619 186379 172622
rect 411253 172546 411319 172549
rect 409860 172544 411319 172546
rect 409860 172488 411258 172544
rect 411314 172488 411319 172544
rect 409860 172486 411319 172488
rect 411253 172483 411319 172486
rect 189398 171602 190072 171662
rect 186313 171594 186379 171597
rect 189398 171594 189458 171602
rect 186313 171592 189458 171594
rect 186313 171536 186318 171592
rect 186374 171536 189458 171592
rect 186313 171534 189458 171536
rect 186313 171531 186379 171534
rect 411253 170506 411319 170509
rect 409860 170504 411319 170506
rect 409860 170448 411258 170504
rect 411314 170448 411319 170504
rect 409860 170446 411319 170448
rect 411253 170443 411319 170446
rect 189398 170378 190072 170438
rect 186313 170370 186379 170373
rect 189398 170370 189458 170378
rect 186313 170368 189458 170370
rect 186313 170312 186318 170368
rect 186374 170312 189458 170368
rect 186313 170310 189458 170312
rect 186313 170307 186379 170310
rect 189398 169290 190072 169350
rect 186313 169282 186379 169285
rect 189398 169282 189458 169290
rect 186313 169280 189458 169282
rect 186313 169224 186318 169280
rect 186374 169224 189458 169280
rect 186313 169222 189458 169224
rect 186313 169219 186379 169222
rect 411253 168602 411319 168605
rect 409860 168600 411319 168602
rect 409860 168544 411258 168600
rect 411314 168544 411319 168600
rect 409860 168542 411319 168544
rect 411253 168539 411319 168542
rect 189398 168202 190072 168262
rect 186405 168194 186471 168197
rect 189398 168194 189458 168202
rect 186405 168192 189458 168194
rect 186405 168136 186410 168192
rect 186466 168136 189458 168192
rect 186405 168134 189458 168136
rect 186405 168131 186471 168134
rect 186313 167106 186379 167109
rect 186313 167104 189642 167106
rect 186313 167048 186318 167104
rect 186374 167078 189642 167104
rect 186374 167048 190164 167078
rect 186313 167046 190164 167048
rect 186313 167043 186379 167046
rect 189582 167018 190164 167046
rect 411253 166562 411319 166565
rect 409860 166560 411319 166562
rect 409860 166504 411258 166560
rect 411314 166504 411319 166560
rect 409860 166502 411319 166504
rect 411253 166499 411319 166502
rect 189398 165890 190072 165950
rect 186313 165882 186379 165885
rect 189398 165882 189458 165890
rect 186313 165880 189458 165882
rect 186313 165824 186318 165880
rect 186374 165824 189458 165880
rect 186313 165822 189458 165824
rect 186313 165819 186379 165822
rect 583520 165732 584960 165972
rect 189398 164802 190072 164862
rect 186313 164794 186379 164797
rect 189398 164794 189458 164802
rect 186313 164792 189458 164794
rect 186313 164736 186318 164792
rect 186374 164736 189458 164792
rect 186313 164734 189458 164736
rect 186313 164731 186379 164734
rect 411253 164658 411319 164661
rect 409860 164656 411319 164658
rect 409860 164600 411258 164656
rect 411314 164600 411319 164656
rect 409860 164598 411319 164600
rect 411253 164595 411319 164598
rect 189398 163714 190072 163774
rect 186313 163706 186379 163709
rect 189398 163706 189458 163714
rect 186313 163704 189458 163706
rect 186313 163648 186318 163704
rect 186374 163648 189458 163704
rect 186313 163646 189458 163648
rect 186313 163643 186379 163646
rect -960 162740 480 162980
rect 411253 162618 411319 162621
rect 409860 162616 411319 162618
rect 409860 162560 411258 162616
rect 411314 162560 411319 162616
rect 409860 162558 411319 162560
rect 411253 162555 411319 162558
rect 189398 162490 190072 162550
rect 186405 162482 186471 162485
rect 189398 162482 189458 162490
rect 186405 162480 189458 162482
rect 186405 162424 186410 162480
rect 186466 162424 189458 162480
rect 186405 162422 189458 162424
rect 186405 162419 186471 162422
rect 186313 161530 186379 161533
rect 186313 161528 189642 161530
rect 186313 161472 186318 161528
rect 186374 161502 189642 161528
rect 186374 161472 190164 161502
rect 186313 161470 190164 161472
rect 186313 161467 186379 161470
rect 189582 161442 190164 161470
rect 411253 160714 411319 160717
rect 409860 160712 411319 160714
rect 409860 160656 411258 160712
rect 411314 160656 411319 160712
rect 409860 160654 411319 160656
rect 411253 160651 411319 160654
rect 189398 160314 190072 160374
rect 186313 160306 186379 160309
rect 189398 160306 189458 160314
rect 186313 160304 189458 160306
rect 186313 160248 186318 160304
rect 186374 160248 189458 160304
rect 186313 160246 189458 160248
rect 186313 160243 186379 160246
rect 189398 159090 190072 159150
rect 186313 159082 186379 159085
rect 189398 159082 189458 159090
rect 186313 159080 189458 159082
rect 186313 159024 186318 159080
rect 186374 159024 189458 159080
rect 186313 159022 189458 159024
rect 186313 159019 186379 159022
rect 411253 158810 411319 158813
rect 409860 158808 411319 158810
rect 409860 158752 411258 158808
rect 411314 158752 411319 158808
rect 409860 158750 411319 158752
rect 411253 158747 411319 158750
rect 189398 158002 190072 158062
rect 186313 157994 186379 157997
rect 189398 157994 189458 158002
rect 186313 157992 189458 157994
rect 186313 157936 186318 157992
rect 186374 157936 189458 157992
rect 186313 157934 189458 157936
rect 186313 157931 186379 157934
rect 189398 156914 190072 156974
rect 186313 156906 186379 156909
rect 189398 156906 189458 156914
rect 186313 156904 189458 156906
rect 186313 156848 186318 156904
rect 186374 156848 189458 156904
rect 186313 156846 189458 156848
rect 186313 156843 186379 156846
rect 411253 156770 411319 156773
rect 409860 156768 411319 156770
rect 409860 156712 411258 156768
rect 411314 156712 411319 156768
rect 409860 156710 411319 156712
rect 411253 156707 411319 156710
rect 189398 155826 190072 155886
rect 186405 155818 186471 155821
rect 189398 155818 189458 155826
rect 186405 155816 189458 155818
rect 186405 155760 186410 155816
rect 186466 155760 189458 155816
rect 186405 155758 189458 155760
rect 186405 155755 186471 155758
rect 411253 154866 411319 154869
rect 409860 154864 411319 154866
rect 409860 154808 411258 154864
rect 411314 154808 411319 154864
rect 409860 154806 411319 154808
rect 411253 154803 411319 154806
rect 186313 154730 186379 154733
rect 186313 154728 189642 154730
rect 186313 154672 186318 154728
rect 186374 154702 189642 154728
rect 186374 154672 190164 154702
rect 186313 154670 190164 154672
rect 186313 154667 186379 154670
rect 189582 154642 190164 154670
rect 189398 153514 190072 153574
rect 186313 153506 186379 153509
rect 189398 153506 189458 153514
rect 186313 153504 189458 153506
rect 186313 153448 186318 153504
rect 186374 153448 189458 153504
rect 186313 153446 189458 153448
rect 186313 153443 186379 153446
rect 411253 152826 411319 152829
rect 409860 152824 411319 152826
rect 409860 152768 411258 152824
rect 411314 152768 411319 152824
rect 409860 152766 411319 152768
rect 411253 152763 411319 152766
rect 580349 152690 580415 152693
rect 583520 152690 584960 152780
rect 580349 152688 584960 152690
rect 580349 152632 580354 152688
rect 580410 152632 584960 152688
rect 580349 152630 584960 152632
rect 580349 152627 580415 152630
rect 583520 152540 584960 152630
rect 189398 152426 190072 152486
rect 186313 152418 186379 152421
rect 189398 152418 189458 152426
rect 186313 152416 189458 152418
rect 186313 152360 186318 152416
rect 186374 152360 189458 152416
rect 186313 152358 189458 152360
rect 186313 152355 186379 152358
rect 189398 151202 190072 151262
rect 186313 151194 186379 151197
rect 189398 151194 189458 151202
rect 186313 151192 189458 151194
rect 186313 151136 186318 151192
rect 186374 151136 189458 151192
rect 186313 151134 189458 151136
rect 186313 151131 186379 151134
rect 411253 150922 411319 150925
rect 409860 150920 411319 150922
rect 409860 150864 411258 150920
rect 411314 150864 411319 150920
rect 409860 150862 411319 150864
rect 411253 150859 411319 150862
rect 189398 150114 190072 150174
rect 186405 150106 186471 150109
rect 189398 150106 189458 150114
rect 186405 150104 189458 150106
rect 186405 150048 186410 150104
rect 186466 150048 189458 150104
rect 186405 150046 189458 150048
rect 186405 150043 186471 150046
rect -960 149684 480 149924
rect 186313 149154 186379 149157
rect 186313 149152 189642 149154
rect 186313 149096 186318 149152
rect 186374 149126 189642 149152
rect 186374 149096 190164 149126
rect 186313 149094 190164 149096
rect 186313 149091 186379 149094
rect 189582 149066 190164 149094
rect 411253 148882 411319 148885
rect 409860 148880 411319 148882
rect 409860 148824 411258 148880
rect 411314 148824 411319 148880
rect 409860 148822 411319 148824
rect 411253 148819 411319 148822
rect 189398 147802 190072 147862
rect 186313 147794 186379 147797
rect 189398 147794 189458 147802
rect 186313 147792 189458 147794
rect 186313 147736 186318 147792
rect 186374 147736 189458 147792
rect 186313 147734 189458 147736
rect 186313 147731 186379 147734
rect 411253 146978 411319 146981
rect 409860 146976 411319 146978
rect 409860 146920 411258 146976
rect 411314 146920 411319 146976
rect 409860 146918 411319 146920
rect 411253 146915 411319 146918
rect 189398 146714 190072 146774
rect 186313 146706 186379 146709
rect 189398 146706 189458 146714
rect 186313 146704 189458 146706
rect 186313 146648 186318 146704
rect 186374 146648 189458 146704
rect 186313 146646 189458 146648
rect 186313 146643 186379 146646
rect 189398 145626 190072 145686
rect 186313 145618 186379 145621
rect 189398 145618 189458 145626
rect 186313 145616 189458 145618
rect 186313 145560 186318 145616
rect 186374 145560 189458 145616
rect 186313 145558 189458 145560
rect 186313 145555 186379 145558
rect 411253 144938 411319 144941
rect 409860 144936 411319 144938
rect 409860 144880 411258 144936
rect 411314 144880 411319 144936
rect 409860 144878 411319 144880
rect 411253 144875 411319 144878
rect 189398 144538 190072 144598
rect 186313 144530 186379 144533
rect 189398 144530 189458 144538
rect 186313 144528 189458 144530
rect 186313 144472 186318 144528
rect 186374 144472 189458 144528
rect 186313 144470 189458 144472
rect 186313 144467 186379 144470
rect 189398 143314 190072 143374
rect 186405 143306 186471 143309
rect 189398 143306 189458 143314
rect 186405 143304 189458 143306
rect 186405 143248 186410 143304
rect 186466 143248 189458 143304
rect 186405 143246 189458 143248
rect 186405 143243 186471 143246
rect 411253 143034 411319 143037
rect 409860 143032 411319 143034
rect 409860 142976 411258 143032
rect 411314 142976 411319 143032
rect 409860 142974 411319 142976
rect 411253 142971 411319 142974
rect 189398 142226 190072 142286
rect 186313 142218 186379 142221
rect 189398 142218 189458 142226
rect 186313 142216 189458 142218
rect 186313 142160 186318 142216
rect 186374 142160 189458 142216
rect 186313 142158 189458 142160
rect 186313 142155 186379 142158
rect 189398 141138 190072 141198
rect 187325 141130 187391 141133
rect 189398 141130 189458 141138
rect 411253 141130 411319 141133
rect 187325 141128 189458 141130
rect 187325 141072 187330 141128
rect 187386 141072 189458 141128
rect 187325 141070 189458 141072
rect 409860 141128 411319 141130
rect 409860 141072 411258 141128
rect 411314 141072 411319 141128
rect 409860 141070 411319 141072
rect 187325 141067 187391 141070
rect 411253 141067 411319 141070
rect 189398 139914 190072 139974
rect 186313 139906 186379 139909
rect 189398 139906 189458 139914
rect 186313 139904 189458 139906
rect 186313 139848 186318 139904
rect 186374 139848 189458 139904
rect 186313 139846 189458 139848
rect 186313 139843 186379 139846
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 411253 139090 411319 139093
rect 409860 139088 411319 139090
rect 409860 139032 411258 139088
rect 411314 139032 411319 139088
rect 409860 139030 411319 139032
rect 411253 139027 411319 139030
rect 189398 138826 190072 138886
rect 186313 138818 186379 138821
rect 189398 138818 189458 138826
rect 186313 138816 189458 138818
rect 186313 138760 186318 138816
rect 186374 138760 189458 138816
rect 186313 138758 189458 138760
rect 186313 138755 186379 138758
rect 189398 137738 190072 137798
rect 186313 137730 186379 137733
rect 189398 137730 189458 137738
rect 186313 137728 189458 137730
rect 186313 137672 186318 137728
rect 186374 137672 189458 137728
rect 186313 137670 189458 137672
rect 186313 137667 186379 137670
rect 411253 137186 411319 137189
rect 409860 137184 411319 137186
rect 409860 137128 411258 137184
rect 411314 137128 411319 137184
rect 409860 137126 411319 137128
rect 411253 137123 411319 137126
rect -960 136628 480 136868
rect 189398 136514 190072 136574
rect 186405 136506 186471 136509
rect 189398 136506 189458 136514
rect 186405 136504 189458 136506
rect 186405 136448 186410 136504
rect 186466 136448 189458 136504
rect 186405 136446 189458 136448
rect 186405 136443 186471 136446
rect 189398 135426 190072 135486
rect 186313 135418 186379 135421
rect 189398 135418 189458 135426
rect 186313 135416 189458 135418
rect 186313 135360 186318 135416
rect 186374 135360 189458 135416
rect 186313 135358 189458 135360
rect 186313 135355 186379 135358
rect 411253 135146 411319 135149
rect 409860 135144 411319 135146
rect 409860 135088 411258 135144
rect 411314 135088 411319 135144
rect 409860 135086 411319 135088
rect 411253 135083 411319 135086
rect 189398 134338 190072 134398
rect 186313 134330 186379 134333
rect 189398 134330 189458 134338
rect 186313 134328 189458 134330
rect 186313 134272 186318 134328
rect 186374 134272 189458 134328
rect 186313 134270 189458 134272
rect 186313 134267 186379 134270
rect 189398 133250 190072 133310
rect 186313 133242 186379 133245
rect 189398 133242 189458 133250
rect 411253 133242 411319 133245
rect 186313 133240 189458 133242
rect 186313 133184 186318 133240
rect 186374 133184 189458 133240
rect 186313 133182 189458 133184
rect 409860 133240 411319 133242
rect 409860 133184 411258 133240
rect 411314 133184 411319 133240
rect 409860 133182 411319 133184
rect 186313 133179 186379 133182
rect 411253 133179 411319 133182
rect 189398 132026 190072 132086
rect 186313 132018 186379 132021
rect 189398 132018 189458 132026
rect 186313 132016 189458 132018
rect 186313 131960 186318 132016
rect 186374 131960 189458 132016
rect 186313 131958 189458 131960
rect 186313 131955 186379 131958
rect 412173 131202 412239 131205
rect 409860 131200 412239 131202
rect 409860 131144 412178 131200
rect 412234 131144 412239 131200
rect 409860 131142 412239 131144
rect 412173 131139 412239 131142
rect 189398 130938 190072 130998
rect 187417 130930 187483 130933
rect 189398 130930 189458 130938
rect 187417 130928 189458 130930
rect 187417 130872 187422 130928
rect 187478 130872 189458 130928
rect 187417 130870 189458 130872
rect 187417 130867 187483 130870
rect 189398 129850 190072 129910
rect 186313 129842 186379 129845
rect 189398 129842 189458 129850
rect 129598 129782 130210 129842
rect 129598 129676 129658 129782
rect 130150 129706 130210 129782
rect 186313 129840 189458 129842
rect 186313 129784 186318 129840
rect 186374 129784 189458 129840
rect 186313 129782 189458 129784
rect 186313 129779 186379 129782
rect 131113 129706 131179 129709
rect 130150 129704 131179 129706
rect 130150 129648 131118 129704
rect 131174 129648 131179 129704
rect 130150 129646 131179 129648
rect 131113 129643 131179 129646
rect 411253 129298 411319 129301
rect 409860 129296 411319 129298
rect 409860 129240 411258 129296
rect 411314 129240 411319 129296
rect 409860 129238 411319 129240
rect 411253 129235 411319 129238
rect 131849 129162 131915 129165
rect 130518 129160 131915 129162
rect 130518 129134 131854 129160
rect 129904 129104 131854 129134
rect 131910 129104 131915 129160
rect 129904 129102 131915 129104
rect 129904 129074 130578 129102
rect 131849 129099 131915 129102
rect 437473 128754 437539 128757
rect 440006 128754 440066 129132
rect 437473 128752 440066 128754
rect 437473 128696 437478 128752
rect 437534 128696 440066 128752
rect 437473 128694 440066 128696
rect 437473 128691 437539 128694
rect 189398 128626 190072 128686
rect 131205 128618 131271 128621
rect 130518 128616 131271 128618
rect 130518 128590 131210 128616
rect 129904 128560 131210 128590
rect 131266 128560 131271 128616
rect 129904 128558 131271 128560
rect 129904 128530 130578 128558
rect 131205 128555 131271 128558
rect 186313 128618 186379 128621
rect 189398 128618 189458 128626
rect 186313 128616 189458 128618
rect 186313 128560 186318 128616
rect 186374 128560 189458 128616
rect 186313 128558 189458 128560
rect 186313 128555 186379 128558
rect 131757 127938 131823 127941
rect 130518 127936 131823 127938
rect 130518 127910 131762 127936
rect 129904 127880 131762 127910
rect 131818 127880 131823 127936
rect 129904 127878 131823 127880
rect 129904 127850 130578 127878
rect 131757 127875 131823 127878
rect 189398 127538 190072 127598
rect 186313 127530 186379 127533
rect 189398 127530 189458 127538
rect 186313 127528 189458 127530
rect 186313 127472 186318 127528
rect 186374 127472 189458 127528
rect 186313 127470 189458 127472
rect 186313 127467 186379 127470
rect 131205 127394 131271 127397
rect 130518 127392 131271 127394
rect 130518 127366 131210 127392
rect 129904 127336 131210 127366
rect 131266 127336 131271 127392
rect 129904 127334 131271 127336
rect 129904 127306 130578 127334
rect 131205 127331 131271 127334
rect 437473 127394 437539 127397
rect 440006 127394 440066 127636
rect 437473 127392 440066 127394
rect 437473 127336 437478 127392
rect 437534 127336 440066 127392
rect 437473 127334 440066 127336
rect 437473 127331 437539 127334
rect 411253 127258 411319 127261
rect 409860 127256 411319 127258
rect 409860 127200 411258 127256
rect 411314 127200 411319 127256
rect 409860 127198 411319 127200
rect 411253 127195 411319 127198
rect 131205 126850 131271 126853
rect 130518 126848 131271 126850
rect 130518 126822 131210 126848
rect 129904 126792 131210 126822
rect 131266 126792 131271 126848
rect 129904 126790 131271 126792
rect 129904 126762 130578 126790
rect 131205 126787 131271 126790
rect 189398 126450 190072 126510
rect 186313 126442 186379 126445
rect 189398 126442 189458 126450
rect 186313 126440 189458 126442
rect 186313 126384 186318 126440
rect 186374 126384 189458 126440
rect 186313 126382 189458 126384
rect 186313 126379 186379 126382
rect 131113 126170 131179 126173
rect 130518 126168 131179 126170
rect 130518 126142 131118 126168
rect 129904 126112 131118 126142
rect 131174 126112 131179 126168
rect 129904 126110 131179 126112
rect 129904 126082 130578 126110
rect 131113 126107 131179 126110
rect 539317 126034 539383 126037
rect 580349 126034 580415 126037
rect 583520 126034 584960 126124
rect 539317 126032 539426 126034
rect 437473 125898 437539 125901
rect 440006 125898 440066 126004
rect 539317 125976 539322 126032
rect 539378 125976 539426 126032
rect 539317 125971 539426 125976
rect 580349 126032 584960 126034
rect 580349 125976 580354 126032
rect 580410 125976 584960 126032
rect 580349 125974 584960 125976
rect 580349 125971 580415 125974
rect 437473 125896 440066 125898
rect 437473 125840 437478 125896
rect 437534 125840 440066 125896
rect 437473 125838 440066 125840
rect 437473 125835 437539 125838
rect 131113 125626 131179 125629
rect 130150 125624 131179 125626
rect 130150 125598 131118 125624
rect 129966 125592 131118 125598
rect 129904 125568 131118 125592
rect 131174 125568 131179 125624
rect 129904 125566 131179 125568
rect 129904 125538 130210 125566
rect 131113 125563 131179 125566
rect 129904 125532 130026 125538
rect 539366 125460 539426 125971
rect 583520 125884 584960 125974
rect 411253 125354 411319 125357
rect 409860 125352 411319 125354
rect 409860 125296 411258 125352
rect 411314 125296 411319 125352
rect 409860 125294 411319 125296
rect 411253 125291 411319 125294
rect 189398 125226 190072 125286
rect 186313 125218 186379 125221
rect 189398 125218 189458 125226
rect 186313 125216 189458 125218
rect 186313 125160 186318 125216
rect 186374 125160 189458 125216
rect 186313 125158 189458 125160
rect 186313 125155 186379 125158
rect 131573 125082 131639 125085
rect 130518 125080 131639 125082
rect 130518 125054 131578 125080
rect 129904 125024 131578 125054
rect 131634 125024 131639 125080
rect 129904 125022 131639 125024
rect 129904 124994 130578 125022
rect 131573 125019 131639 125022
rect 131205 124538 131271 124541
rect 130518 124536 131271 124538
rect 130518 124510 131210 124536
rect 129904 124480 131210 124510
rect 131266 124480 131271 124536
rect 129904 124478 131271 124480
rect 129904 124450 130578 124478
rect 131205 124475 131271 124478
rect 187509 124266 187575 124269
rect 437473 124266 437539 124269
rect 440006 124266 440066 124508
rect 187509 124264 189642 124266
rect 187509 124208 187514 124264
rect 187570 124238 189642 124264
rect 437473 124264 440066 124266
rect 187570 124208 190164 124238
rect 187509 124206 190164 124208
rect 187509 124203 187575 124206
rect 189582 124178 190164 124206
rect 437473 124208 437478 124264
rect 437534 124208 440066 124264
rect 437473 124206 440066 124208
rect 437473 124203 437539 124206
rect 131757 123858 131823 123861
rect 130518 123856 131823 123858
rect 130518 123830 131762 123856
rect -960 123572 480 123812
rect 129904 123800 131762 123830
rect 131818 123800 131823 123856
rect 129904 123798 131823 123800
rect 129904 123770 130578 123798
rect 131757 123795 131823 123798
rect 131113 123314 131179 123317
rect 411253 123314 411319 123317
rect 130518 123312 131179 123314
rect 130518 123286 131118 123312
rect 129904 123256 131118 123286
rect 131174 123256 131179 123312
rect 129904 123254 131179 123256
rect 409860 123312 411319 123314
rect 409860 123256 411258 123312
rect 411314 123256 411319 123312
rect 409860 123254 411319 123256
rect 129904 123226 130578 123254
rect 131113 123251 131179 123254
rect 411253 123251 411319 123254
rect 189398 123050 190072 123110
rect 186313 123042 186379 123045
rect 189398 123042 189458 123050
rect 186313 123040 189458 123042
rect 186313 122984 186318 123040
rect 186374 122984 189458 123040
rect 186313 122982 189458 122984
rect 437473 123042 437539 123045
rect 437473 123040 440066 123042
rect 437473 122984 437478 123040
rect 437534 122984 440066 123040
rect 437473 122982 440066 122984
rect 186313 122979 186379 122982
rect 437473 122979 437539 122982
rect 440006 122876 440066 122982
rect 131205 122770 131271 122773
rect 130518 122768 131271 122770
rect 130518 122742 131210 122768
rect 129904 122712 131210 122742
rect 131266 122712 131271 122768
rect 129904 122710 131271 122712
rect 129904 122682 130578 122710
rect 131205 122707 131271 122710
rect 131481 122090 131547 122093
rect 130518 122088 131547 122090
rect 130518 122062 131486 122088
rect 129904 122032 131486 122062
rect 131542 122032 131547 122088
rect 129904 122030 131547 122032
rect 129904 122002 130578 122030
rect 131481 122027 131547 122030
rect 189398 121962 190072 122022
rect 186313 121954 186379 121957
rect 189398 121954 189458 121962
rect 186313 121952 189458 121954
rect 186313 121896 186318 121952
rect 186374 121896 189458 121952
rect 186313 121894 189458 121896
rect 186313 121891 186379 121894
rect 131113 121546 131179 121549
rect 130518 121544 131179 121546
rect 130518 121518 131118 121544
rect 129904 121488 131118 121518
rect 131174 121488 131179 121544
rect 129904 121486 131179 121488
rect 129904 121458 130578 121486
rect 131113 121483 131179 121486
rect 411253 121410 411319 121413
rect 409860 121408 411319 121410
rect 409860 121352 411258 121408
rect 411314 121352 411319 121408
rect 409860 121350 411319 121352
rect 411253 121347 411319 121350
rect 131205 121002 131271 121005
rect 130518 121000 131271 121002
rect 130518 120974 131210 121000
rect 129904 120944 131210 120974
rect 131266 120944 131271 121000
rect 129904 120942 131271 120944
rect 129904 120914 130578 120942
rect 131205 120939 131271 120942
rect 438485 120866 438551 120869
rect 440006 120866 440066 121380
rect 438485 120864 440066 120866
rect 438485 120808 438490 120864
rect 438546 120808 440066 120864
rect 438485 120806 440066 120808
rect 438485 120803 438551 120806
rect 189398 120738 190072 120798
rect 186957 120730 187023 120733
rect 189398 120730 189458 120738
rect 186957 120728 189458 120730
rect 186957 120672 186962 120728
rect 187018 120672 189458 120728
rect 186957 120670 189458 120672
rect 186957 120667 187023 120670
rect 131113 120322 131179 120325
rect 130518 120320 131179 120322
rect 130518 120294 131118 120320
rect 129904 120264 131118 120294
rect 131174 120264 131179 120320
rect 129904 120262 131179 120264
rect 129904 120234 130578 120262
rect 131113 120259 131179 120262
rect 132309 119778 132375 119781
rect 130518 119776 132375 119778
rect 130518 119750 132314 119776
rect 129904 119720 132314 119750
rect 132370 119720 132375 119776
rect 129904 119718 132375 119720
rect 129904 119690 130578 119718
rect 132309 119715 132375 119718
rect 189398 119650 190072 119710
rect 186313 119642 186379 119645
rect 189398 119642 189458 119650
rect 186313 119640 189458 119642
rect 186313 119584 186318 119640
rect 186374 119584 189458 119640
rect 186313 119582 189458 119584
rect 186313 119579 186379 119582
rect 411253 119506 411319 119509
rect 409860 119504 411319 119506
rect 409860 119448 411258 119504
rect 411314 119448 411319 119504
rect 409860 119446 411319 119448
rect 411253 119443 411319 119446
rect 131113 119234 131179 119237
rect 130518 119232 131179 119234
rect 130518 119206 131118 119232
rect 129904 119176 131118 119206
rect 131174 119176 131179 119232
rect 129904 119174 131179 119176
rect 129904 119146 130578 119174
rect 131113 119171 131179 119174
rect 438393 119234 438459 119237
rect 440006 119234 440066 119748
rect 438393 119232 440066 119234
rect 438393 119176 438398 119232
rect 438454 119176 440066 119232
rect 438393 119174 440066 119176
rect 438393 119171 438459 119174
rect 129968 118562 130578 118622
rect 130518 118554 130578 118562
rect 189398 118562 190072 118622
rect 131205 118554 131271 118557
rect 130518 118552 131271 118554
rect 130518 118496 131210 118552
rect 131266 118496 131271 118552
rect 130518 118494 131271 118496
rect 131205 118491 131271 118494
rect 186405 118554 186471 118557
rect 189398 118554 189458 118562
rect 186405 118552 189458 118554
rect 186405 118496 186410 118552
rect 186466 118496 189458 118552
rect 186405 118494 189458 118496
rect 186405 118491 186471 118494
rect 131297 118010 131363 118013
rect 130518 118008 131363 118010
rect 130518 117982 131302 118008
rect 129904 117952 131302 117982
rect 131358 117952 131363 118008
rect 129904 117950 131363 117952
rect 129904 117922 130578 117950
rect 131297 117947 131363 117950
rect 438301 117738 438367 117741
rect 440006 117738 440066 118252
rect 438301 117736 440066 117738
rect 438301 117680 438306 117736
rect 438362 117680 440066 117736
rect 438301 117678 440066 117680
rect 438301 117675 438367 117678
rect 131113 117466 131179 117469
rect 412265 117466 412331 117469
rect 130518 117464 131179 117466
rect 130518 117438 131118 117464
rect 129904 117408 131118 117438
rect 131174 117408 131179 117464
rect 129904 117406 131179 117408
rect 409860 117464 412331 117466
rect 409860 117408 412270 117464
rect 412326 117408 412331 117464
rect 409860 117406 412331 117408
rect 129904 117378 130578 117406
rect 131113 117403 131179 117406
rect 412265 117403 412331 117406
rect 189398 117338 190072 117398
rect 186313 117330 186379 117333
rect 189398 117330 189458 117338
rect 186313 117328 189458 117330
rect 186313 117272 186318 117328
rect 186374 117272 189458 117328
rect 186313 117270 189458 117272
rect 186313 117267 186379 117270
rect 131205 116922 131271 116925
rect 130518 116920 131271 116922
rect 130518 116894 131210 116920
rect 129904 116864 131210 116894
rect 131266 116864 131271 116920
rect 129904 116862 131271 116864
rect 129904 116834 130578 116862
rect 131205 116859 131271 116862
rect 189398 116250 190072 116310
rect 131113 116242 131179 116245
rect 130518 116240 131179 116242
rect 130518 116214 131118 116240
rect 129904 116184 131118 116214
rect 131174 116184 131179 116240
rect 129904 116182 131179 116184
rect 129904 116154 130578 116182
rect 131113 116179 131179 116182
rect 186313 116242 186379 116245
rect 189398 116242 189458 116250
rect 186313 116240 189458 116242
rect 186313 116184 186318 116240
rect 186374 116184 189458 116240
rect 186313 116182 189458 116184
rect 186313 116179 186379 116182
rect 438209 116106 438275 116109
rect 440006 116106 440066 116620
rect 542445 116378 542511 116381
rect 539948 116376 542511 116378
rect 539948 116320 542450 116376
rect 542506 116320 542511 116376
rect 539948 116318 542511 116320
rect 542445 116315 542511 116318
rect 438209 116104 440066 116106
rect 438209 116048 438214 116104
rect 438270 116048 440066 116104
rect 438209 116046 440066 116048
rect 438209 116043 438275 116046
rect 132309 115698 132375 115701
rect 130518 115696 132375 115698
rect 130518 115670 132314 115696
rect 129904 115640 132314 115670
rect 132370 115640 132375 115696
rect 129904 115638 132375 115640
rect 129904 115610 130578 115638
rect 132309 115635 132375 115638
rect 411253 115562 411319 115565
rect 409860 115560 411319 115562
rect 409860 115504 411258 115560
rect 411314 115504 411319 115560
rect 409860 115502 411319 115504
rect 411253 115499 411319 115502
rect 189398 115162 190072 115222
rect 131205 115154 131271 115157
rect 130518 115152 131271 115154
rect 130518 115126 131210 115152
rect 129904 115096 131210 115126
rect 131266 115096 131271 115152
rect 129904 115094 131271 115096
rect 129904 115066 130578 115094
rect 131205 115091 131271 115094
rect 186313 115154 186379 115157
rect 189398 115154 189458 115162
rect 186313 115152 189458 115154
rect 186313 115096 186318 115152
rect 186374 115096 189458 115152
rect 186313 115094 189458 115096
rect 186313 115091 186379 115094
rect 438117 114610 438183 114613
rect 440006 114610 440066 115124
rect 438117 114608 440066 114610
rect 438117 114552 438122 114608
rect 438178 114552 440066 114608
rect 438117 114550 440066 114552
rect 438117 114547 438183 114550
rect 131205 114474 131271 114477
rect 130518 114472 131271 114474
rect 130518 114446 131210 114472
rect 129904 114416 131210 114446
rect 131266 114416 131271 114472
rect 129904 114414 131271 114416
rect 129904 114386 130578 114414
rect 131205 114411 131271 114414
rect 189398 114074 190072 114134
rect 186313 114066 186379 114069
rect 189398 114066 189458 114074
rect 186313 114064 189458 114066
rect 186313 114008 186318 114064
rect 186374 114008 189458 114064
rect 186313 114006 189458 114008
rect 437473 114066 437539 114069
rect 437473 114064 440066 114066
rect 437473 114008 437478 114064
rect 437534 114008 440066 114064
rect 437473 114006 440066 114008
rect 186313 114003 186379 114006
rect 437473 114003 437539 114006
rect 131113 113930 131179 113933
rect 130518 113928 131179 113930
rect 130518 113902 131118 113928
rect 129904 113872 131118 113902
rect 131174 113872 131179 113928
rect 129904 113870 131179 113872
rect 129904 113842 130578 113870
rect 131113 113867 131179 113870
rect 411253 113522 411319 113525
rect 409860 113520 411319 113522
rect 409860 113464 411258 113520
rect 411314 113464 411319 113520
rect 440006 113492 440066 114006
rect 409860 113462 411319 113464
rect 411253 113459 411319 113462
rect 131297 113386 131363 113389
rect 130518 113384 131363 113386
rect 130518 113358 131302 113384
rect 129904 113328 131302 113358
rect 131358 113328 131363 113384
rect 129904 113326 131363 113328
rect 129904 113298 130578 113326
rect 131297 113323 131363 113326
rect 189398 112850 190072 112910
rect 131205 112842 131271 112845
rect 130518 112840 131271 112842
rect 130518 112814 131210 112840
rect 129904 112784 131210 112814
rect 131266 112784 131271 112840
rect 129904 112782 131271 112784
rect 129904 112754 130578 112782
rect 131205 112779 131271 112782
rect 186405 112842 186471 112845
rect 189398 112842 189458 112850
rect 186405 112840 189458 112842
rect 186405 112784 186410 112840
rect 186466 112784 189458 112840
rect 186405 112782 189458 112784
rect 580257 112842 580323 112845
rect 583520 112842 584960 112932
rect 580257 112840 584960 112842
rect 580257 112784 580262 112840
rect 580318 112784 584960 112840
rect 580257 112782 584960 112784
rect 186405 112779 186471 112782
rect 580257 112779 580323 112782
rect 583520 112692 584960 112782
rect 437473 112570 437539 112573
rect 437473 112568 440066 112570
rect 437473 112512 437478 112568
rect 437534 112512 440066 112568
rect 437473 112510 440066 112512
rect 437473 112507 437539 112510
rect 131113 112162 131179 112165
rect 130518 112160 131179 112162
rect 130518 112134 131118 112160
rect 129904 112104 131118 112134
rect 131174 112104 131179 112160
rect 129904 112102 131179 112104
rect 129904 112074 130578 112102
rect 131113 112099 131179 112102
rect 440006 111996 440066 112510
rect 186313 111890 186379 111893
rect 186313 111888 189642 111890
rect 186313 111832 186318 111888
rect 186374 111862 189642 111888
rect 186374 111832 190164 111862
rect 186313 111830 190164 111832
rect 186313 111827 186379 111830
rect 189582 111802 190164 111830
rect 131205 111618 131271 111621
rect 411897 111618 411963 111621
rect 130518 111616 131271 111618
rect 130518 111590 131210 111616
rect 129904 111560 131210 111590
rect 131266 111560 131271 111616
rect 129904 111558 131271 111560
rect 409860 111616 411963 111618
rect 409860 111560 411902 111616
rect 411958 111560 411963 111616
rect 409860 111558 411963 111560
rect 129904 111530 130578 111558
rect 131205 111555 131271 111558
rect 411897 111555 411963 111558
rect 131113 111074 131179 111077
rect 130518 111072 131179 111074
rect 130518 111046 131118 111072
rect 129904 111016 131118 111046
rect 131174 111016 131179 111072
rect 129904 111014 131179 111016
rect 129904 110986 130578 111014
rect 131113 111011 131179 111014
rect -960 110516 480 110756
rect 189398 110674 190072 110734
rect 187049 110666 187115 110669
rect 189398 110666 189458 110674
rect 187049 110664 189458 110666
rect 187049 110608 187054 110664
rect 187110 110608 189458 110664
rect 187049 110606 189458 110608
rect 187049 110603 187115 110606
rect 131205 110394 131271 110397
rect 130518 110392 131271 110394
rect 130518 110366 131210 110392
rect 129904 110336 131210 110366
rect 131266 110336 131271 110392
rect 129904 110334 131271 110336
rect 129904 110306 130578 110334
rect 131205 110331 131271 110334
rect 437473 110258 437539 110261
rect 440006 110258 440066 110364
rect 437473 110256 440066 110258
rect 437473 110200 437478 110256
rect 437534 110200 440066 110256
rect 437473 110198 440066 110200
rect 437473 110195 437539 110198
rect 131205 109850 131271 109853
rect 130518 109848 131271 109850
rect 130518 109822 131210 109848
rect 129904 109792 131210 109822
rect 131266 109792 131271 109848
rect 129904 109790 131271 109792
rect 129904 109762 130578 109790
rect 131205 109787 131271 109790
rect 411253 109578 411319 109581
rect 409860 109576 411319 109578
rect 409860 109520 411258 109576
rect 411314 109520 411319 109576
rect 409860 109518 411319 109520
rect 411253 109515 411319 109518
rect 189398 109450 190072 109510
rect 186313 109442 186379 109445
rect 189398 109442 189458 109450
rect 186313 109440 189458 109442
rect 186313 109384 186318 109440
rect 186374 109384 189458 109440
rect 186313 109382 189458 109384
rect 186313 109379 186379 109382
rect 131113 109306 131179 109309
rect 130518 109304 131179 109306
rect 130518 109278 131118 109304
rect 129904 109248 131118 109278
rect 131174 109248 131179 109304
rect 129904 109246 131179 109248
rect 129904 109218 130578 109246
rect 131113 109243 131179 109246
rect 437473 109034 437539 109037
rect 437473 109032 440066 109034
rect 437473 108976 437478 109032
rect 437534 108976 440066 109032
rect 437473 108974 440066 108976
rect 437473 108971 437539 108974
rect 440006 108868 440066 108974
rect 131205 108626 131271 108629
rect 130518 108624 131271 108626
rect 130518 108598 131210 108624
rect 129904 108568 131210 108598
rect 131266 108568 131271 108624
rect 129904 108566 131271 108568
rect 129904 108538 130578 108566
rect 131205 108563 131271 108566
rect 189398 108362 190072 108422
rect 186313 108354 186379 108357
rect 189398 108354 189458 108362
rect 186313 108352 189458 108354
rect 186313 108296 186318 108352
rect 186374 108296 189458 108352
rect 186313 108294 189458 108296
rect 186313 108291 186379 108294
rect 131113 108082 131179 108085
rect 130518 108080 131179 108082
rect 130518 108054 131118 108080
rect 129904 108024 131118 108054
rect 131174 108024 131179 108080
rect 129904 108022 131179 108024
rect 129904 107994 130578 108022
rect 131113 108019 131179 108022
rect 411253 107674 411319 107677
rect 409860 107672 411319 107674
rect 409860 107616 411258 107672
rect 411314 107616 411319 107672
rect 409860 107614 411319 107616
rect 411253 107611 411319 107614
rect 131205 107538 131271 107541
rect 130518 107536 131271 107538
rect 130518 107510 131210 107536
rect 129904 107480 131210 107510
rect 131266 107480 131271 107536
rect 129904 107478 131271 107480
rect 129904 107450 130578 107478
rect 131205 107475 131271 107478
rect 437473 107402 437539 107405
rect 437473 107400 440066 107402
rect 437473 107344 437478 107400
rect 437534 107344 440066 107400
rect 437473 107342 440066 107344
rect 437473 107339 437539 107342
rect 189398 107274 190072 107334
rect 186313 107266 186379 107269
rect 189398 107266 189458 107274
rect 186313 107264 189458 107266
rect 186313 107208 186318 107264
rect 186374 107208 189458 107264
rect 440006 107236 440066 107342
rect 542353 107266 542419 107269
rect 539948 107264 542419 107266
rect 186313 107206 189458 107208
rect 539948 107208 542358 107264
rect 542414 107208 542419 107264
rect 539948 107206 542419 107208
rect 186313 107203 186379 107206
rect 542353 107203 542419 107206
rect 131113 106994 131179 106997
rect 130518 106992 131179 106994
rect 130518 106966 131118 106992
rect 129904 106936 131118 106966
rect 131174 106936 131179 106992
rect 129904 106934 131179 106936
rect 129904 106906 130578 106934
rect 131113 106931 131179 106934
rect 131297 106314 131363 106317
rect 130150 106312 131363 106314
rect 130150 106280 131302 106312
rect 129904 106256 131302 106280
rect 131358 106256 131363 106312
rect 129904 106254 131363 106256
rect 129904 106220 130210 106254
rect 131297 106251 131363 106254
rect 436737 106178 436803 106181
rect 436737 106176 440066 106178
rect 436737 106120 436742 106176
rect 436798 106120 440066 106176
rect 436737 106118 440066 106120
rect 436737 106115 436803 106118
rect 189398 106050 190072 106110
rect 186405 106042 186471 106045
rect 189398 106042 189458 106050
rect 186405 106040 189458 106042
rect 186405 105984 186410 106040
rect 186466 105984 189458 106040
rect 186405 105982 189458 105984
rect 186405 105979 186471 105982
rect 131205 105770 131271 105773
rect 130518 105768 131271 105770
rect 130518 105742 131210 105768
rect 129904 105712 131210 105742
rect 131266 105712 131271 105768
rect 440006 105740 440066 106118
rect 129904 105710 131271 105712
rect 129904 105682 130578 105710
rect 131205 105707 131271 105710
rect 411989 105634 412055 105637
rect 409860 105632 412055 105634
rect 409860 105576 411994 105632
rect 412050 105576 412055 105632
rect 409860 105574 412055 105576
rect 411989 105571 412055 105574
rect 131113 105226 131179 105229
rect 130518 105224 131179 105226
rect 130518 105198 131118 105224
rect 129904 105168 131118 105198
rect 131174 105168 131179 105224
rect 129904 105166 131179 105168
rect 129904 105138 130578 105166
rect 131113 105163 131179 105166
rect 189398 104962 190072 105022
rect 186313 104954 186379 104957
rect 189398 104954 189458 104962
rect 186313 104952 189458 104954
rect 186313 104896 186318 104952
rect 186374 104896 189458 104952
rect 186313 104894 189458 104896
rect 186313 104891 186379 104894
rect 131205 104546 131271 104549
rect 130518 104544 131271 104546
rect 130518 104518 131210 104544
rect 129904 104488 131210 104518
rect 131266 104488 131271 104544
rect 129904 104486 131271 104488
rect 129904 104458 130578 104486
rect 131205 104483 131271 104486
rect 437473 104546 437539 104549
rect 437473 104544 440066 104546
rect 437473 104488 437478 104544
rect 437534 104488 440066 104544
rect 437473 104486 440066 104488
rect 437473 104483 437539 104486
rect 440006 104108 440066 104486
rect 131113 104002 131179 104005
rect 130518 104000 131179 104002
rect 130518 103974 131118 104000
rect 129904 103944 131118 103974
rect 131174 103944 131179 104000
rect 129904 103942 131179 103944
rect 129904 103914 130578 103942
rect 131113 103939 131179 103942
rect 189398 103874 190072 103934
rect 187141 103866 187207 103869
rect 189398 103866 189458 103874
rect 187141 103864 189458 103866
rect 187141 103808 187146 103864
rect 187202 103808 189458 103864
rect 187141 103806 189458 103808
rect 187141 103803 187207 103806
rect 411253 103730 411319 103733
rect 409860 103728 411319 103730
rect 409860 103672 411258 103728
rect 411314 103672 411319 103728
rect 409860 103670 411319 103672
rect 411253 103667 411319 103670
rect 131205 103458 131271 103461
rect 130518 103456 131271 103458
rect 130518 103430 131210 103456
rect 129904 103400 131210 103430
rect 131266 103400 131271 103456
rect 129904 103398 131271 103400
rect 129904 103370 130578 103398
rect 131205 103395 131271 103398
rect 437657 103050 437723 103053
rect 437657 103048 440066 103050
rect 437657 102992 437662 103048
rect 437718 102992 440066 103048
rect 437657 102990 440066 102992
rect 437657 102987 437723 102990
rect 189398 102786 190072 102846
rect 131389 102778 131455 102781
rect 130518 102776 131455 102778
rect 130518 102750 131394 102776
rect 129904 102720 131394 102750
rect 131450 102720 131455 102776
rect 129904 102718 131455 102720
rect 129904 102690 130578 102718
rect 131389 102715 131455 102718
rect 186313 102778 186379 102781
rect 189398 102778 189458 102786
rect 186313 102776 189458 102778
rect 186313 102720 186318 102776
rect 186374 102720 189458 102776
rect 186313 102718 189458 102720
rect 186313 102715 186379 102718
rect 440006 102612 440066 102990
rect 131113 102234 131179 102237
rect 130518 102232 131179 102234
rect 130518 102206 131118 102232
rect 129904 102176 131118 102206
rect 131174 102176 131179 102232
rect 129904 102174 131179 102176
rect 129904 102146 130578 102174
rect 131113 102171 131179 102174
rect 411253 101826 411319 101829
rect 409860 101824 411319 101826
rect 409860 101768 411258 101824
rect 411314 101768 411319 101824
rect 409860 101766 411319 101768
rect 411253 101763 411319 101766
rect 131941 101690 132007 101693
rect 130518 101688 132007 101690
rect 130518 101662 131946 101688
rect 129904 101632 131946 101662
rect 132002 101632 132007 101688
rect 129904 101630 132007 101632
rect 129904 101602 130578 101630
rect 131941 101627 132007 101630
rect 189398 101562 190072 101622
rect 186313 101554 186379 101557
rect 189398 101554 189458 101562
rect 186313 101552 189458 101554
rect 186313 101496 186318 101552
rect 186374 101496 189458 101552
rect 186313 101494 189458 101496
rect 437473 101554 437539 101557
rect 437473 101552 440066 101554
rect 437473 101496 437478 101552
rect 437534 101496 440066 101552
rect 437473 101494 440066 101496
rect 186313 101491 186379 101494
rect 437473 101491 437539 101494
rect 131205 101146 131271 101149
rect 130518 101144 131271 101146
rect 130518 101118 131210 101144
rect 129904 101088 131210 101118
rect 131266 101088 131271 101144
rect 129904 101086 131271 101088
rect 129904 101058 130578 101086
rect 131205 101083 131271 101086
rect 440006 100980 440066 101494
rect 189398 100474 190072 100534
rect 131205 100466 131271 100469
rect 130518 100464 131271 100466
rect 130518 100438 131210 100464
rect 129904 100408 131210 100438
rect 131266 100408 131271 100464
rect 129904 100406 131271 100408
rect 129904 100378 130578 100406
rect 131205 100403 131271 100406
rect 186405 100466 186471 100469
rect 189398 100466 189458 100474
rect 186405 100464 189458 100466
rect 186405 100408 186410 100464
rect 186466 100408 189458 100464
rect 186405 100406 189458 100408
rect 186405 100403 186471 100406
rect 437473 100058 437539 100061
rect 437473 100056 440066 100058
rect 437473 100000 437478 100056
rect 437534 100000 440066 100056
rect 437473 99998 440066 100000
rect 437473 99995 437539 99998
rect 131113 99922 131179 99925
rect 130518 99920 131179 99922
rect 130518 99894 131118 99920
rect 129904 99864 131118 99894
rect 131174 99864 131179 99920
rect 129904 99862 131179 99864
rect 129904 99834 130578 99862
rect 131113 99859 131179 99862
rect 412081 99786 412147 99789
rect 409860 99784 412147 99786
rect 409860 99728 412086 99784
rect 412142 99728 412147 99784
rect 409860 99726 412147 99728
rect 412081 99723 412147 99726
rect 186313 99514 186379 99517
rect 186313 99512 189642 99514
rect 186313 99456 186318 99512
rect 186374 99486 189642 99512
rect 186374 99456 190164 99486
rect 440006 99484 440066 99998
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 186313 99454 190164 99456
rect 186313 99451 186379 99454
rect 189582 99426 190164 99454
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 131665 99378 131731 99381
rect 130518 99376 131731 99378
rect 130518 99350 131670 99376
rect 129904 99320 131670 99350
rect 131726 99320 131731 99376
rect 583520 99364 584960 99454
rect 129904 99318 131731 99320
rect 129904 99290 130578 99318
rect 131665 99315 131731 99318
rect 131205 98698 131271 98701
rect 130518 98696 131271 98698
rect 130518 98670 131210 98696
rect 129904 98640 131210 98670
rect 131266 98640 131271 98696
rect 129904 98638 131271 98640
rect 129904 98610 130578 98638
rect 131205 98635 131271 98638
rect 189398 98162 190072 98222
rect 131113 98154 131179 98157
rect 130518 98152 131179 98154
rect 130518 98126 131118 98152
rect 129904 98096 131118 98126
rect 131174 98096 131179 98152
rect 129904 98094 131179 98096
rect 129904 98066 130578 98094
rect 131113 98091 131179 98094
rect 186313 98154 186379 98157
rect 189398 98154 189458 98162
rect 542353 98154 542419 98157
rect 186313 98152 189458 98154
rect 186313 98096 186318 98152
rect 186374 98096 189458 98152
rect 186313 98094 189458 98096
rect 539948 98152 542419 98154
rect 539948 98096 542358 98152
rect 542414 98096 542419 98152
rect 539948 98094 542419 98096
rect 186313 98091 186379 98094
rect 542353 98091 542419 98094
rect 412357 97882 412423 97885
rect 409860 97880 412423 97882
rect 409860 97824 412362 97880
rect 412418 97824 412423 97880
rect 409860 97822 412423 97824
rect 412357 97819 412423 97822
rect 437473 97746 437539 97749
rect 440006 97746 440066 97852
rect 437473 97744 440066 97746
rect -960 97460 480 97700
rect 437473 97688 437478 97744
rect 437534 97688 440066 97744
rect 437473 97686 440066 97688
rect 437473 97683 437539 97686
rect 131205 97610 131271 97613
rect 130518 97608 131271 97610
rect 130518 97582 131210 97608
rect 129904 97552 131210 97582
rect 131266 97552 131271 97608
rect 129904 97550 131271 97552
rect 129904 97522 130578 97550
rect 131205 97547 131271 97550
rect 189398 97074 190072 97134
rect 131573 97066 131639 97069
rect 130518 97064 131639 97066
rect 130518 97038 131578 97064
rect 129904 97008 131578 97038
rect 131634 97008 131639 97064
rect 129904 97006 131639 97008
rect 129904 96978 130578 97006
rect 131573 97003 131639 97006
rect 186313 97066 186379 97069
rect 189398 97066 189458 97074
rect 186313 97064 189458 97066
rect 186313 97008 186318 97064
rect 186374 97008 189458 97064
rect 186313 97006 189458 97008
rect 186313 97003 186379 97006
rect 437473 96522 437539 96525
rect 437473 96520 440066 96522
rect 437473 96464 437478 96520
rect 437534 96464 440066 96520
rect 437473 96462 440066 96464
rect 437473 96459 437539 96462
rect 131205 96386 131271 96389
rect 130518 96384 131271 96386
rect 130518 96358 131210 96384
rect 129904 96328 131210 96358
rect 131266 96328 131271 96384
rect 440006 96356 440066 96462
rect 129904 96326 131271 96328
rect 129904 96298 130578 96326
rect 131205 96323 131271 96326
rect 189398 95986 190072 96046
rect 186313 95978 186379 95981
rect 189398 95978 189458 95986
rect 186313 95976 189458 95978
rect 186313 95920 186318 95976
rect 186374 95920 189458 95976
rect 186313 95918 189458 95920
rect 186313 95915 186379 95918
rect 131113 95842 131179 95845
rect 411253 95842 411319 95845
rect 130518 95840 131179 95842
rect 130518 95814 131118 95840
rect 129904 95784 131118 95814
rect 131174 95784 131179 95840
rect 129904 95782 131179 95784
rect 409860 95840 411319 95842
rect 409860 95784 411258 95840
rect 411314 95784 411319 95840
rect 409860 95782 411319 95784
rect 129904 95754 130578 95782
rect 131113 95779 131179 95782
rect 411253 95779 411319 95782
rect 131389 95298 131455 95301
rect 130518 95296 131455 95298
rect 130518 95270 131394 95296
rect 129904 95240 131394 95270
rect 131450 95240 131455 95296
rect 129904 95238 131455 95240
rect 129904 95210 130578 95238
rect 131389 95235 131455 95238
rect 437473 95162 437539 95165
rect 437473 95160 440066 95162
rect 437473 95104 437478 95160
rect 437534 95104 440066 95160
rect 437473 95102 440066 95104
rect 437473 95099 437539 95102
rect 189398 94762 190072 94822
rect 186313 94754 186379 94757
rect 189398 94754 189458 94762
rect 186313 94752 189458 94754
rect 186313 94696 186318 94752
rect 186374 94696 189458 94752
rect 440006 94724 440066 95102
rect 186313 94694 189458 94696
rect 186313 94691 186379 94694
rect 131205 94618 131271 94621
rect 130518 94616 131271 94618
rect 130518 94590 131210 94616
rect 129904 94560 131210 94590
rect 131266 94560 131271 94616
rect 129904 94558 131271 94560
rect 129904 94530 130578 94558
rect 131205 94555 131271 94558
rect 131113 94074 131179 94077
rect 130518 94072 131179 94074
rect 130518 94046 131118 94072
rect 129904 94016 131118 94046
rect 131174 94016 131179 94072
rect 129904 94014 131179 94016
rect 129904 93986 130578 94014
rect 131113 94011 131179 94014
rect 411253 93938 411319 93941
rect 409860 93936 411319 93938
rect 409860 93880 411258 93936
rect 411314 93880 411319 93936
rect 409860 93878 411319 93880
rect 411253 93875 411319 93878
rect 189398 93674 190072 93734
rect 186405 93666 186471 93669
rect 189398 93666 189458 93674
rect 186405 93664 189458 93666
rect 186405 93608 186410 93664
rect 186466 93608 189458 93664
rect 186405 93606 189458 93608
rect 186405 93603 186471 93606
rect 131205 93530 131271 93533
rect 130518 93528 131271 93530
rect 130518 93502 131210 93528
rect 129904 93472 131210 93502
rect 131266 93472 131271 93528
rect 129904 93470 131271 93472
rect 129904 93442 130578 93470
rect 131205 93467 131271 93470
rect 437473 93530 437539 93533
rect 437473 93528 440066 93530
rect 437473 93472 437478 93528
rect 437534 93472 440066 93528
rect 437473 93470 440066 93472
rect 437473 93467 437539 93470
rect 440006 93228 440066 93470
rect 131113 92850 131179 92853
rect 130518 92848 131179 92850
rect 130518 92822 131118 92848
rect 129904 92792 131118 92822
rect 131174 92792 131179 92848
rect 129904 92790 131179 92792
rect 129904 92762 130578 92790
rect 131113 92787 131179 92790
rect 189398 92586 190072 92646
rect 186313 92578 186379 92581
rect 189398 92578 189458 92586
rect 186313 92576 189458 92578
rect 186313 92520 186318 92576
rect 186374 92520 189458 92576
rect 186313 92518 189458 92520
rect 186313 92515 186379 92518
rect 131205 92306 131271 92309
rect 130518 92304 131271 92306
rect 130518 92278 131210 92304
rect 129904 92248 131210 92278
rect 131266 92248 131271 92304
rect 129904 92246 131271 92248
rect 129904 92218 130578 92246
rect 131205 92243 131271 92246
rect 437473 92034 437539 92037
rect 437473 92032 440066 92034
rect 437473 91976 437478 92032
rect 437534 91976 440066 92032
rect 437473 91974 440066 91976
rect 437473 91971 437539 91974
rect 411253 91898 411319 91901
rect 409860 91896 411319 91898
rect 409860 91840 411258 91896
rect 411314 91840 411319 91896
rect 409860 91838 411319 91840
rect 411253 91835 411319 91838
rect 131113 91762 131179 91765
rect 130518 91760 131179 91762
rect 130518 91734 131118 91760
rect 129904 91704 131118 91734
rect 131174 91704 131179 91760
rect 129904 91702 131179 91704
rect 129904 91674 130578 91702
rect 131113 91699 131179 91702
rect 440006 91596 440066 91974
rect 189398 91498 190072 91558
rect 186313 91490 186379 91493
rect 189398 91490 189458 91498
rect 186313 91488 189458 91490
rect 186313 91432 186318 91488
rect 186374 91432 189458 91488
rect 186313 91430 189458 91432
rect 186313 91427 186379 91430
rect 132217 91218 132283 91221
rect 130518 91216 132283 91218
rect 130518 91190 132222 91216
rect 129904 91160 132222 91190
rect 132278 91160 132283 91216
rect 129904 91158 132283 91160
rect 129904 91130 130578 91158
rect 132217 91155 132283 91158
rect 132217 90538 132283 90541
rect 130518 90536 132283 90538
rect 130518 90510 132222 90536
rect 129904 90480 132222 90510
rect 132278 90480 132283 90536
rect 129904 90478 132283 90480
rect 129904 90450 130578 90478
rect 132217 90475 132283 90478
rect 437473 90538 437539 90541
rect 437473 90536 440066 90538
rect 437473 90480 437478 90536
rect 437534 90480 440066 90536
rect 437473 90478 440066 90480
rect 437473 90475 437539 90478
rect 189398 90274 190072 90334
rect 186313 90266 186379 90269
rect 189398 90266 189458 90274
rect 186313 90264 189458 90266
rect 186313 90208 186318 90264
rect 186374 90208 189458 90264
rect 186313 90206 189458 90208
rect 186313 90203 186379 90206
rect 440006 90100 440066 90478
rect 131205 89994 131271 89997
rect 411253 89994 411319 89997
rect 130518 89992 131271 89994
rect 130518 89966 131210 89992
rect 129904 89936 131210 89966
rect 131266 89936 131271 89992
rect 129904 89934 131271 89936
rect 409860 89992 411319 89994
rect 409860 89936 411258 89992
rect 411314 89936 411319 89992
rect 409860 89934 411319 89936
rect 129904 89906 130578 89934
rect 131205 89931 131271 89934
rect 411253 89931 411319 89934
rect 131205 89450 131271 89453
rect 130518 89448 131271 89450
rect 130518 89422 131210 89448
rect 129904 89392 131210 89422
rect 131266 89392 131271 89448
rect 129904 89390 131271 89392
rect 129904 89362 130578 89390
rect 131205 89387 131271 89390
rect 189398 89186 190072 89246
rect 186313 89178 186379 89181
rect 189398 89178 189458 89186
rect 186313 89176 189458 89178
rect 186313 89120 186318 89176
rect 186374 89120 189458 89176
rect 186313 89118 189458 89120
rect 186313 89115 186379 89118
rect 437473 89042 437539 89045
rect 542445 89042 542511 89045
rect 437473 89040 440066 89042
rect 437473 88984 437478 89040
rect 437534 88984 440066 89040
rect 437473 88982 440066 88984
rect 539948 89040 542511 89042
rect 539948 88984 542450 89040
rect 542506 88984 542511 89040
rect 539948 88982 542511 88984
rect 437473 88979 437539 88982
rect 131113 88770 131179 88773
rect 130518 88768 131179 88770
rect 130518 88742 131118 88768
rect 129904 88712 131118 88742
rect 131174 88712 131179 88768
rect 129904 88710 131179 88712
rect 129904 88682 130578 88710
rect 131113 88707 131179 88710
rect 440006 88468 440066 88982
rect 542445 88979 542511 88982
rect 131205 88226 131271 88229
rect 130518 88224 131271 88226
rect 130518 88198 131210 88224
rect 129904 88168 131210 88198
rect 131266 88168 131271 88224
rect 129904 88166 131271 88168
rect 129904 88138 130578 88166
rect 131205 88163 131271 88166
rect 189398 88098 190072 88158
rect 186313 88090 186379 88093
rect 189398 88090 189458 88098
rect 186313 88088 189458 88090
rect 186313 88032 186318 88088
rect 186374 88032 189458 88088
rect 186313 88030 189458 88032
rect 186313 88027 186379 88030
rect 411253 87954 411319 87957
rect 409860 87952 411319 87954
rect 409860 87896 411258 87952
rect 411314 87896 411319 87952
rect 409860 87894 411319 87896
rect 411253 87891 411319 87894
rect 131113 87682 131179 87685
rect 130518 87680 131179 87682
rect 130518 87654 131118 87680
rect 129904 87624 131118 87654
rect 131174 87624 131179 87680
rect 129904 87622 131179 87624
rect 129904 87594 130578 87622
rect 131113 87619 131179 87622
rect 437473 87546 437539 87549
rect 437473 87544 440066 87546
rect 437473 87488 437478 87544
rect 437534 87488 440066 87544
rect 437473 87486 440066 87488
rect 437473 87483 437539 87486
rect 131297 87002 131363 87005
rect 130518 87000 131363 87002
rect 130518 86974 131302 87000
rect 129904 86944 131302 86974
rect 131358 86944 131363 87000
rect 129904 86942 131363 86944
rect 129904 86914 130578 86942
rect 131297 86939 131363 86942
rect 187233 87002 187299 87005
rect 187233 87000 189642 87002
rect 187233 86944 187238 87000
rect 187294 86974 189642 87000
rect 187294 86944 190164 86974
rect 440006 86972 440066 87486
rect 187233 86942 190164 86944
rect 187233 86939 187299 86942
rect 189582 86914 190164 86942
rect 131113 86458 131179 86461
rect 130518 86456 131179 86458
rect 130518 86430 131118 86456
rect 129904 86400 131118 86430
rect 131174 86400 131179 86456
rect 129904 86398 131179 86400
rect 129904 86370 130578 86398
rect 131113 86395 131179 86398
rect 580257 86186 580323 86189
rect 583520 86186 584960 86276
rect 580257 86184 584960 86186
rect 580257 86128 580262 86184
rect 580318 86128 584960 86184
rect 580257 86126 584960 86128
rect 580257 86123 580323 86126
rect 411253 86050 411319 86053
rect 409860 86048 411319 86050
rect 409860 85992 411258 86048
rect 411314 85992 411319 86048
rect 583520 86036 584960 86126
rect 409860 85990 411319 85992
rect 411253 85987 411319 85990
rect 131205 85914 131271 85917
rect 130518 85912 131271 85914
rect 130518 85886 131210 85912
rect 129904 85856 131210 85886
rect 131266 85856 131271 85912
rect 129904 85854 131271 85856
rect 129904 85826 130578 85854
rect 131205 85851 131271 85854
rect 189398 85786 190072 85846
rect 186313 85778 186379 85781
rect 189398 85778 189458 85786
rect 186313 85776 189458 85778
rect 186313 85720 186318 85776
rect 186374 85720 189458 85776
rect 186313 85718 189458 85720
rect 186313 85715 186379 85718
rect 437473 85506 437539 85509
rect 437473 85504 440066 85506
rect 437473 85448 437478 85504
rect 437534 85448 440066 85504
rect 437473 85446 440066 85448
rect 437473 85443 437539 85446
rect 131205 85370 131271 85373
rect 130518 85368 131271 85370
rect 130518 85342 131210 85368
rect 129904 85312 131210 85342
rect 131266 85312 131271 85368
rect 440006 85340 440066 85446
rect 129904 85310 131271 85312
rect 129904 85282 130578 85310
rect 131205 85307 131271 85310
rect -960 84540 480 84780
rect 189398 84698 190072 84758
rect 131113 84690 131179 84693
rect 130518 84688 131179 84690
rect 130518 84662 131118 84688
rect 129904 84632 131118 84662
rect 131174 84632 131179 84688
rect 129904 84630 131179 84632
rect 129904 84602 130578 84630
rect 131113 84627 131179 84630
rect 186313 84690 186379 84693
rect 189398 84690 189458 84698
rect 186313 84688 189458 84690
rect 186313 84632 186318 84688
rect 186374 84632 189458 84688
rect 186313 84630 189458 84632
rect 186313 84627 186379 84630
rect 131205 84146 131271 84149
rect 411253 84146 411319 84149
rect 130518 84144 131271 84146
rect 130518 84118 131210 84144
rect 129904 84088 131210 84118
rect 131266 84088 131271 84144
rect 129904 84086 131271 84088
rect 409860 84144 411319 84146
rect 409860 84088 411258 84144
rect 411314 84088 411319 84144
rect 409860 84086 411319 84088
rect 129904 84058 130578 84086
rect 131205 84083 131271 84086
rect 411253 84083 411319 84086
rect 437473 84146 437539 84149
rect 437473 84144 440066 84146
rect 437473 84088 437478 84144
rect 437534 84088 440066 84144
rect 437473 84086 440066 84088
rect 437473 84083 437539 84086
rect 440006 83844 440066 84086
rect 131573 83602 131639 83605
rect 130518 83600 131639 83602
rect 130518 83574 131578 83600
rect 129904 83544 131578 83574
rect 131634 83544 131639 83600
rect 129904 83542 131639 83544
rect 129904 83514 130578 83542
rect 131573 83539 131639 83542
rect 189398 83474 190072 83534
rect 187325 83466 187391 83469
rect 189398 83466 189458 83474
rect 187325 83464 189458 83466
rect 187325 83408 187330 83464
rect 187386 83408 189458 83464
rect 187325 83406 189458 83408
rect 187325 83403 187391 83406
rect 131113 82922 131179 82925
rect 130518 82920 131179 82922
rect 130518 82894 131118 82920
rect 129904 82864 131118 82894
rect 131174 82864 131179 82920
rect 129904 82862 131179 82864
rect 129904 82834 130578 82862
rect 131113 82859 131179 82862
rect 437473 82514 437539 82517
rect 437473 82512 440066 82514
rect 437473 82456 437478 82512
rect 437534 82456 440066 82512
rect 437473 82454 440066 82456
rect 437473 82451 437539 82454
rect 189398 82386 190072 82446
rect 131205 82378 131271 82381
rect 130518 82376 131271 82378
rect 130518 82350 131210 82376
rect 129904 82320 131210 82350
rect 131266 82320 131271 82376
rect 129904 82318 131271 82320
rect 129904 82290 130578 82318
rect 131205 82315 131271 82318
rect 186313 82378 186379 82381
rect 189398 82378 189458 82386
rect 186313 82376 189458 82378
rect 186313 82320 186318 82376
rect 186374 82320 189458 82376
rect 186313 82318 189458 82320
rect 186313 82315 186379 82318
rect 440006 82212 440066 82454
rect 411253 82106 411319 82109
rect 409860 82104 411319 82106
rect 409860 82048 411258 82104
rect 411314 82048 411319 82104
rect 409860 82046 411319 82048
rect 411253 82043 411319 82046
rect 131113 81834 131179 81837
rect 130518 81832 131179 81834
rect 130518 81806 131118 81832
rect 129904 81776 131118 81806
rect 131174 81776 131179 81832
rect 129904 81774 131179 81776
rect 129904 81746 130578 81774
rect 131113 81771 131179 81774
rect 189398 81298 190072 81358
rect 186313 81290 186379 81293
rect 189398 81290 189458 81298
rect 186313 81288 189458 81290
rect 186313 81232 186318 81288
rect 186374 81232 189458 81288
rect 186313 81230 189458 81232
rect 186313 81227 186379 81230
rect 131205 81154 131271 81157
rect 130518 81152 131271 81154
rect 130518 81126 131210 81152
rect 129904 81096 131210 81126
rect 131266 81096 131271 81152
rect 129904 81094 131271 81096
rect 129904 81066 130578 81094
rect 131205 81091 131271 81094
rect 437473 81018 437539 81021
rect 437473 81016 440066 81018
rect 437473 80960 437478 81016
rect 437534 80960 440066 81016
rect 437473 80958 440066 80960
rect 437473 80955 437539 80958
rect 440006 80716 440066 80958
rect 131113 80610 131179 80613
rect 130518 80608 131179 80610
rect 130518 80582 131118 80608
rect 129904 80552 131118 80582
rect 131174 80552 131179 80608
rect 129904 80550 131179 80552
rect 129904 80522 130578 80550
rect 131113 80547 131179 80550
rect 189398 80210 190072 80270
rect 187417 80202 187483 80205
rect 189398 80202 189458 80210
rect 412541 80202 412607 80205
rect 187417 80200 189458 80202
rect 187417 80144 187422 80200
rect 187478 80144 189458 80200
rect 187417 80142 189458 80144
rect 409860 80200 412607 80202
rect 409860 80144 412546 80200
rect 412602 80144 412607 80200
rect 409860 80142 412607 80144
rect 187417 80139 187483 80142
rect 412541 80139 412607 80142
rect 542537 80066 542603 80069
rect 539948 80064 542603 80066
rect 539948 80008 542542 80064
rect 542598 80008 542603 80064
rect 539948 80006 542603 80008
rect 542537 80003 542603 80006
rect 129968 79938 130578 79998
rect 130518 79930 130578 79938
rect 131205 79930 131271 79933
rect 130518 79928 131271 79930
rect 130518 79872 131210 79928
rect 131266 79872 131271 79928
rect 130518 79870 131271 79872
rect 131205 79867 131271 79870
rect 437473 79658 437539 79661
rect 437473 79656 440066 79658
rect 437473 79600 437478 79656
rect 437534 79600 440066 79656
rect 437473 79598 440066 79600
rect 437473 79595 437539 79598
rect 131113 79522 131179 79525
rect 130518 79520 131179 79522
rect 130518 79494 131118 79520
rect 129904 79464 131118 79494
rect 131174 79464 131179 79520
rect 129904 79462 131179 79464
rect 129904 79434 130578 79462
rect 131113 79459 131179 79462
rect 440006 79220 440066 79598
rect 189398 78986 190072 79046
rect 186313 78978 186379 78981
rect 189398 78978 189458 78986
rect 186313 78976 189458 78978
rect 186313 78920 186318 78976
rect 186374 78920 189458 78976
rect 186313 78918 189458 78920
rect 186313 78915 186379 78918
rect 131297 78842 131363 78845
rect 130518 78840 131363 78842
rect 130518 78814 131302 78840
rect 129904 78784 131302 78814
rect 131358 78784 131363 78840
rect 129904 78782 131363 78784
rect 129904 78754 130578 78782
rect 131297 78779 131363 78782
rect 131205 78298 131271 78301
rect 130518 78296 131271 78298
rect 130518 78270 131210 78296
rect 129904 78240 131210 78270
rect 131266 78240 131271 78296
rect 129904 78238 131271 78240
rect 129904 78210 130578 78238
rect 131205 78235 131271 78238
rect 411253 78162 411319 78165
rect 409860 78160 411319 78162
rect 409860 78104 411258 78160
rect 411314 78104 411319 78160
rect 409860 78102 411319 78104
rect 411253 78099 411319 78102
rect 437473 78162 437539 78165
rect 437473 78160 440066 78162
rect 437473 78104 437478 78160
rect 437534 78104 440066 78160
rect 437473 78102 440066 78104
rect 437473 78099 437539 78102
rect 189398 77898 190072 77958
rect 186313 77890 186379 77893
rect 189398 77890 189458 77898
rect 186313 77888 189458 77890
rect 186313 77832 186318 77888
rect 186374 77832 189458 77888
rect 186313 77830 189458 77832
rect 186313 77827 186379 77830
rect 131113 77754 131179 77757
rect 130518 77752 131179 77754
rect 130518 77726 131118 77752
rect 129904 77696 131118 77726
rect 131174 77696 131179 77752
rect 129904 77694 131179 77696
rect 129904 77666 130578 77694
rect 131113 77691 131179 77694
rect 440006 77588 440066 78102
rect 131205 77074 131271 77077
rect 130518 77072 131271 77074
rect 130518 77046 131210 77072
rect 129904 77016 131210 77046
rect 131266 77016 131271 77072
rect 129904 77014 131271 77016
rect 129904 76986 130578 77014
rect 131205 77011 131271 77014
rect 189398 76810 190072 76870
rect 187509 76802 187575 76805
rect 189398 76802 189458 76810
rect 187509 76800 189458 76802
rect 187509 76744 187514 76800
rect 187570 76744 189458 76800
rect 187509 76742 189458 76744
rect 187509 76739 187575 76742
rect 437473 76666 437539 76669
rect 437473 76664 440066 76666
rect 437473 76608 437478 76664
rect 437534 76608 440066 76664
rect 437473 76606 440066 76608
rect 437473 76603 437539 76606
rect 131297 76530 131363 76533
rect 130518 76528 131363 76530
rect 130518 76502 131302 76528
rect 129904 76472 131302 76502
rect 131358 76472 131363 76528
rect 129904 76470 131363 76472
rect 129904 76442 130578 76470
rect 131297 76467 131363 76470
rect 411253 76258 411319 76261
rect 409860 76256 411319 76258
rect 409860 76200 411258 76256
rect 411314 76200 411319 76256
rect 409860 76198 411319 76200
rect 411253 76195 411319 76198
rect 440006 76092 440066 76606
rect 131665 75986 131731 75989
rect 130518 75984 131731 75986
rect 130518 75958 131670 75984
rect 129904 75928 131670 75958
rect 131726 75928 131731 75984
rect 129904 75926 131731 75928
rect 129904 75898 130578 75926
rect 131665 75923 131731 75926
rect 189398 75586 190072 75646
rect 186405 75578 186471 75581
rect 189398 75578 189458 75586
rect 186405 75576 189458 75578
rect 186405 75520 186410 75576
rect 186466 75520 189458 75576
rect 186405 75518 189458 75520
rect 186405 75515 186471 75518
rect 131849 75306 131915 75309
rect 130518 75304 131915 75306
rect 130518 75278 131854 75304
rect 129904 75248 131854 75278
rect 131910 75248 131915 75304
rect 129904 75246 131915 75248
rect 129904 75218 130578 75246
rect 131849 75243 131915 75246
rect 131205 74762 131271 74765
rect 130518 74760 131271 74762
rect 130518 74734 131210 74760
rect 129904 74704 131210 74734
rect 131266 74704 131271 74760
rect 129904 74702 131271 74704
rect 129904 74674 130578 74702
rect 131205 74699 131271 74702
rect 186313 74626 186379 74629
rect 186313 74624 189642 74626
rect 186313 74568 186318 74624
rect 186374 74598 189642 74624
rect 186374 74568 190164 74598
rect 186313 74566 190164 74568
rect 186313 74563 186379 74566
rect 189582 74538 190164 74566
rect 437473 74354 437539 74357
rect 440006 74354 440066 74460
rect 437473 74352 440066 74354
rect 437473 74296 437478 74352
rect 437534 74296 440066 74352
rect 437473 74294 440066 74296
rect 437473 74291 437539 74294
rect 131849 74218 131915 74221
rect 411253 74218 411319 74221
rect 130518 74216 131915 74218
rect 130518 74190 131854 74216
rect 129904 74160 131854 74190
rect 131910 74160 131915 74216
rect 129904 74158 131915 74160
rect 409860 74216 411319 74218
rect 409860 74160 411258 74216
rect 411314 74160 411319 74216
rect 409860 74158 411319 74160
rect 129904 74130 130578 74158
rect 131849 74155 131915 74158
rect 411253 74155 411319 74158
rect 132309 73674 132375 73677
rect 130518 73672 132375 73674
rect 130518 73646 132314 73672
rect 129904 73616 132314 73646
rect 132370 73616 132375 73672
rect 129904 73614 132375 73616
rect 129904 73586 130578 73614
rect 132309 73611 132375 73614
rect 189398 73410 190072 73470
rect 186957 73402 187023 73405
rect 189398 73402 189458 73410
rect 186957 73400 189458 73402
rect 186957 73344 186962 73400
rect 187018 73344 189458 73400
rect 186957 73342 189458 73344
rect 186957 73339 187023 73342
rect 437473 73130 437539 73133
rect 437473 73128 440066 73130
rect 437473 73072 437478 73128
rect 437534 73072 440066 73128
rect 437473 73070 440066 73072
rect 437473 73067 437539 73070
rect 131205 72994 131271 72997
rect 130518 72992 131271 72994
rect 130518 72966 131210 72992
rect 129904 72936 131210 72966
rect 131266 72936 131271 72992
rect 440006 72964 440066 73070
rect 580441 72994 580507 72997
rect 583520 72994 584960 73084
rect 580441 72992 584960 72994
rect 129904 72934 131271 72936
rect 129904 72906 130578 72934
rect 131205 72931 131271 72934
rect 580441 72936 580446 72992
rect 580502 72936 584960 72992
rect 580441 72934 584960 72936
rect 580441 72931 580507 72934
rect 583520 72844 584960 72934
rect 131113 72450 131179 72453
rect 130518 72448 131179 72450
rect 130518 72422 131118 72448
rect 129904 72392 131118 72422
rect 131174 72392 131179 72448
rect 129904 72390 131179 72392
rect 129904 72362 130578 72390
rect 131113 72387 131179 72390
rect 189398 72322 190072 72382
rect 186313 72314 186379 72317
rect 189398 72314 189458 72322
rect 411253 72314 411319 72317
rect 186313 72312 189458 72314
rect 186313 72256 186318 72312
rect 186374 72256 189458 72312
rect 186313 72254 189458 72256
rect 409860 72312 411319 72314
rect 409860 72256 411258 72312
rect 411314 72256 411319 72312
rect 409860 72254 411319 72256
rect 186313 72251 186379 72254
rect 411253 72251 411319 72254
rect 131297 71906 131363 71909
rect 130518 71904 131363 71906
rect 130518 71878 131302 71904
rect 129904 71848 131302 71878
rect 131358 71848 131363 71904
rect 129904 71846 131363 71848
rect 129904 71818 130578 71846
rect 131297 71843 131363 71846
rect -960 71484 480 71724
rect 437473 71498 437539 71501
rect 437473 71496 440066 71498
rect 437473 71440 437478 71496
rect 437534 71440 440066 71496
rect 437473 71438 440066 71440
rect 437473 71435 437539 71438
rect 440006 71332 440066 71438
rect 131205 71226 131271 71229
rect 130518 71224 131271 71226
rect 130518 71198 131210 71224
rect 129904 71168 131210 71198
rect 131266 71168 131271 71224
rect 129904 71166 131271 71168
rect 129904 71138 130578 71166
rect 131205 71163 131271 71166
rect 189398 71098 190072 71158
rect 186313 71090 186379 71093
rect 189398 71090 189458 71098
rect 186313 71088 189458 71090
rect 186313 71032 186318 71088
rect 186374 71032 189458 71088
rect 186313 71030 189458 71032
rect 186313 71027 186379 71030
rect 542629 70954 542695 70957
rect 539948 70952 542695 70954
rect 539948 70896 542634 70952
rect 542690 70896 542695 70952
rect 539948 70894 542695 70896
rect 542629 70891 542695 70894
rect 131113 70682 131179 70685
rect 130518 70680 131179 70682
rect 130518 70654 131118 70680
rect 129904 70624 131118 70654
rect 131174 70624 131179 70680
rect 129904 70622 131179 70624
rect 129904 70594 130578 70622
rect 131113 70619 131179 70622
rect 411345 70274 411411 70277
rect 409860 70272 411411 70274
rect 409860 70216 411350 70272
rect 411406 70216 411411 70272
rect 409860 70214 411411 70216
rect 411345 70211 411411 70214
rect 437473 70274 437539 70277
rect 437473 70272 440066 70274
rect 437473 70216 437478 70272
rect 437534 70216 440066 70272
rect 437473 70214 440066 70216
rect 437473 70211 437539 70214
rect 131205 70138 131271 70141
rect 130518 70136 131271 70138
rect 130518 70110 131210 70136
rect 129904 70080 131210 70110
rect 131266 70080 131271 70136
rect 129904 70078 131271 70080
rect 129904 70050 130578 70078
rect 131205 70075 131271 70078
rect 189398 70010 190072 70070
rect 186313 70002 186379 70005
rect 189398 70002 189458 70010
rect 186313 70000 189458 70002
rect 186313 69944 186318 70000
rect 186374 69944 189458 70000
rect 186313 69942 189458 69944
rect 186313 69939 186379 69942
rect 440006 69836 440066 70214
rect 131113 69458 131179 69461
rect 130518 69456 131179 69458
rect 130518 69430 131118 69456
rect 129904 69400 131118 69430
rect 131174 69400 131179 69456
rect 129904 69398 131179 69400
rect 129904 69370 130578 69398
rect 131113 69395 131179 69398
rect 186405 69050 186471 69053
rect 186405 69048 189826 69050
rect 186405 68992 186410 69048
rect 186466 69022 189826 69048
rect 186466 68992 190010 69022
rect 186405 68990 190010 68992
rect 186405 68987 186471 68990
rect 189766 68982 190010 68990
rect 189766 68962 190072 68982
rect 189950 68922 190072 68962
rect 131205 68914 131271 68917
rect 130518 68912 131271 68914
rect 130518 68886 131210 68912
rect 129904 68856 131210 68886
rect 131266 68856 131271 68912
rect 129904 68854 131271 68856
rect 129904 68826 130578 68854
rect 131205 68851 131271 68854
rect 437473 68642 437539 68645
rect 437473 68640 440066 68642
rect 437473 68584 437478 68640
rect 437534 68584 440066 68640
rect 437473 68582 440066 68584
rect 437473 68579 437539 68582
rect 131389 68370 131455 68373
rect 411253 68370 411319 68373
rect 130518 68368 131455 68370
rect 130518 68342 131394 68368
rect 129904 68312 131394 68342
rect 131450 68312 131455 68368
rect 129904 68310 131455 68312
rect 409860 68368 411319 68370
rect 409860 68312 411258 68368
rect 411314 68312 411319 68368
rect 409860 68310 411319 68312
rect 129904 68282 130578 68310
rect 131389 68307 131455 68310
rect 411253 68307 411319 68310
rect 440006 68204 440066 68582
rect 131113 67826 131179 67829
rect 130518 67824 131179 67826
rect 130518 67798 131118 67824
rect 129904 67768 131118 67798
rect 131174 67768 131179 67824
rect 129904 67766 131179 67768
rect 129904 67738 130578 67766
rect 131113 67763 131179 67766
rect 189398 67698 190072 67758
rect 186313 67690 186379 67693
rect 189398 67690 189458 67698
rect 186313 67688 189458 67690
rect 186313 67632 186318 67688
rect 186374 67632 189458 67688
rect 186313 67630 189458 67632
rect 186313 67627 186379 67630
rect 131205 67146 131271 67149
rect 130518 67144 131271 67146
rect 130518 67118 131210 67144
rect 129904 67088 131210 67118
rect 131266 67088 131271 67144
rect 129904 67086 131271 67088
rect 129904 67058 130578 67086
rect 131205 67083 131271 67086
rect 437473 67146 437539 67149
rect 437473 67144 440066 67146
rect 437473 67088 437478 67144
rect 437534 67088 440066 67144
rect 437473 67086 440066 67088
rect 437473 67083 437539 67086
rect 440006 66708 440066 67086
rect 189398 66610 190072 66670
rect 131113 66602 131179 66605
rect 130518 66600 131179 66602
rect 130518 66574 131118 66600
rect 129904 66544 131118 66574
rect 131174 66544 131179 66600
rect 129904 66542 131179 66544
rect 129904 66514 130578 66542
rect 131113 66539 131179 66542
rect 186313 66602 186379 66605
rect 189398 66602 189458 66610
rect 186313 66600 189458 66602
rect 186313 66544 186318 66600
rect 186374 66544 189458 66600
rect 186313 66542 189458 66544
rect 186313 66539 186379 66542
rect 411253 66466 411319 66469
rect 409860 66464 411319 66466
rect 409860 66408 411258 66464
rect 411314 66408 411319 66464
rect 409860 66406 411319 66408
rect 411253 66403 411319 66406
rect 131205 66058 131271 66061
rect 130518 66056 131271 66058
rect 130518 66030 131210 66056
rect 129904 66000 131210 66030
rect 131266 66000 131271 66056
rect 129904 65998 131271 66000
rect 129904 65970 130578 65998
rect 131205 65995 131271 65998
rect 437473 65650 437539 65653
rect 437473 65648 440066 65650
rect 437473 65592 437478 65648
rect 437534 65592 440066 65648
rect 437473 65590 440066 65592
rect 437473 65587 437539 65590
rect 189398 65522 190072 65582
rect 186313 65514 186379 65517
rect 189398 65514 189458 65522
rect 186313 65512 189458 65514
rect 186313 65456 186318 65512
rect 186374 65456 189458 65512
rect 186313 65454 189458 65456
rect 186313 65451 186379 65454
rect 131113 65378 131179 65381
rect 130518 65376 131179 65378
rect 130518 65350 131118 65376
rect 129904 65320 131118 65350
rect 131174 65320 131179 65376
rect 129904 65318 131179 65320
rect 129904 65290 130578 65318
rect 131113 65315 131179 65318
rect 440006 65076 440066 65590
rect 131205 64834 131271 64837
rect 130518 64832 131271 64834
rect 130518 64806 131210 64832
rect 129904 64776 131210 64806
rect 131266 64776 131271 64832
rect 129904 64774 131271 64776
rect 129904 64746 130578 64774
rect 131205 64771 131271 64774
rect 411253 64426 411319 64429
rect 409860 64424 411319 64426
rect 409860 64368 411258 64424
rect 411314 64368 411319 64424
rect 409860 64366 411319 64368
rect 411253 64363 411319 64366
rect 189398 64298 190072 64358
rect 131297 64290 131363 64293
rect 130518 64288 131363 64290
rect 130518 64262 131302 64288
rect 129904 64232 131302 64262
rect 131358 64232 131363 64288
rect 129904 64230 131363 64232
rect 129904 64202 130578 64230
rect 131297 64227 131363 64230
rect 186313 64290 186379 64293
rect 189398 64290 189458 64298
rect 186313 64288 189458 64290
rect 186313 64232 186318 64288
rect 186374 64232 189458 64288
rect 186313 64230 189458 64232
rect 186313 64227 186379 64230
rect 437473 64154 437539 64157
rect 437473 64152 440066 64154
rect 437473 64096 437478 64152
rect 437534 64096 440066 64152
rect 437473 64094 440066 64096
rect 437473 64091 437539 64094
rect 131113 63746 131179 63749
rect 130518 63744 131179 63746
rect 130518 63718 131118 63744
rect 129904 63688 131118 63718
rect 131174 63688 131179 63744
rect 129904 63686 131179 63688
rect 129904 63658 130578 63686
rect 131113 63683 131179 63686
rect 440006 63580 440066 64094
rect 189398 63210 190072 63270
rect 187141 63202 187207 63205
rect 189398 63202 189458 63210
rect 187141 63200 189458 63202
rect 187141 63144 187146 63200
rect 187202 63144 189458 63200
rect 187141 63142 189458 63144
rect 187141 63139 187207 63142
rect 131205 63066 131271 63069
rect 130518 63064 131271 63066
rect 130518 63038 131210 63064
rect 129904 63008 131210 63038
rect 131266 63008 131271 63064
rect 129904 63006 131271 63008
rect 129904 62978 130578 63006
rect 131205 63003 131271 63006
rect 131941 62522 132007 62525
rect 411253 62522 411319 62525
rect 130518 62520 132007 62522
rect 130518 62494 131946 62520
rect 129904 62464 131946 62494
rect 132002 62464 132007 62520
rect 129904 62462 132007 62464
rect 409860 62520 411319 62522
rect 409860 62464 411258 62520
rect 411314 62464 411319 62520
rect 409860 62462 411319 62464
rect 129904 62434 130578 62462
rect 131941 62459 132007 62462
rect 411253 62459 411319 62462
rect 186313 62250 186379 62253
rect 186313 62248 189642 62250
rect 186313 62192 186318 62248
rect 186374 62222 189642 62248
rect 186374 62192 190164 62222
rect 186313 62190 190164 62192
rect 186313 62187 186379 62190
rect 189582 62162 190164 62190
rect 437473 62114 437539 62117
rect 437473 62112 440066 62114
rect 437473 62056 437478 62112
rect 437534 62056 440066 62112
rect 437473 62054 440066 62056
rect 437473 62051 437539 62054
rect 131205 61978 131271 61981
rect 130518 61976 131271 61978
rect 130518 61950 131210 61976
rect 129904 61920 131210 61950
rect 131266 61920 131271 61976
rect 440006 61948 440066 62054
rect 129904 61918 131271 61920
rect 129904 61890 130578 61918
rect 131205 61915 131271 61918
rect 542721 61842 542787 61845
rect 539948 61840 542787 61842
rect 539948 61784 542726 61840
rect 542782 61784 542787 61840
rect 539948 61782 542787 61784
rect 542721 61779 542787 61782
rect 131113 61298 131179 61301
rect 130518 61296 131179 61298
rect 130518 61270 131118 61296
rect 129904 61240 131118 61270
rect 131174 61240 131179 61296
rect 129904 61238 131179 61240
rect 129904 61210 130578 61238
rect 131113 61235 131179 61238
rect 189398 61034 190072 61094
rect 186313 61026 186379 61029
rect 189398 61026 189458 61034
rect 186313 61024 189458 61026
rect 186313 60968 186318 61024
rect 186374 60968 189458 61024
rect 186313 60966 189458 60968
rect 186313 60963 186379 60966
rect 132033 60754 132099 60757
rect 130150 60752 132099 60754
rect 130150 60720 132038 60752
rect 129904 60696 132038 60720
rect 132094 60696 132099 60752
rect 129904 60694 132099 60696
rect 129904 60660 130210 60694
rect 132033 60691 132099 60694
rect 437473 60618 437539 60621
rect 437473 60616 440066 60618
rect 437473 60560 437478 60616
rect 437534 60560 440066 60616
rect 437473 60558 440066 60560
rect 437473 60555 437539 60558
rect 411253 60482 411319 60485
rect 409860 60480 411319 60482
rect 409860 60424 411258 60480
rect 411314 60424 411319 60480
rect 440006 60452 440066 60558
rect 409860 60422 411319 60424
rect 411253 60419 411319 60422
rect 131205 60210 131271 60213
rect 130518 60208 131271 60210
rect 130518 60182 131210 60208
rect 129904 60152 131210 60182
rect 131266 60152 131271 60208
rect 129904 60150 131271 60152
rect 129904 60122 130578 60150
rect 131205 60147 131271 60150
rect 189398 59810 190072 59870
rect 187049 59802 187115 59805
rect 189398 59802 189458 59810
rect 187049 59800 189458 59802
rect 187049 59744 187054 59800
rect 187110 59744 189458 59800
rect 187049 59742 189458 59744
rect 187049 59739 187115 59742
rect 579797 59666 579863 59669
rect 583520 59666 584960 59756
rect 579797 59664 584960 59666
rect 579797 59608 579802 59664
rect 579858 59608 584960 59664
rect 579797 59606 584960 59608
rect 579797 59603 579863 59606
rect 131113 59530 131179 59533
rect 130518 59528 131179 59530
rect 130518 59502 131118 59528
rect 129904 59472 131118 59502
rect 131174 59472 131179 59528
rect 583520 59516 584960 59606
rect 129904 59470 131179 59472
rect 129904 59442 130578 59470
rect 131113 59467 131179 59470
rect 437473 59258 437539 59261
rect 437473 59256 440066 59258
rect 437473 59200 437478 59256
rect 437534 59200 440066 59256
rect 437473 59198 440066 59200
rect 437473 59195 437539 59198
rect 131573 58986 131639 58989
rect 130518 58984 131639 58986
rect 130518 58958 131578 58984
rect 129904 58928 131578 58958
rect 131634 58928 131639 58984
rect 129904 58926 131639 58928
rect 129904 58898 130578 58926
rect 131573 58923 131639 58926
rect 440006 58820 440066 59198
rect 189398 58722 190072 58782
rect 186313 58714 186379 58717
rect 189398 58714 189458 58722
rect 186313 58712 189458 58714
rect -960 58428 480 58668
rect 186313 58656 186318 58712
rect 186374 58656 189458 58712
rect 186313 58654 189458 58656
rect 186313 58651 186379 58654
rect 411253 58578 411319 58581
rect 409860 58576 411319 58578
rect 409860 58520 411258 58576
rect 411314 58520 411319 58576
rect 409860 58518 411319 58520
rect 411253 58515 411319 58518
rect 131205 58442 131271 58445
rect 130518 58440 131271 58442
rect 130518 58414 131210 58440
rect 129904 58384 131210 58414
rect 131266 58384 131271 58440
rect 129904 58382 131271 58384
rect 129904 58354 130578 58382
rect 131205 58379 131271 58382
rect 131205 57898 131271 57901
rect 130518 57896 131271 57898
rect 130518 57870 131210 57896
rect 129904 57840 131210 57870
rect 131266 57840 131271 57896
rect 129904 57838 131271 57840
rect 129904 57810 130578 57838
rect 131205 57835 131271 57838
rect 189398 57634 190072 57694
rect 186313 57626 186379 57629
rect 189398 57626 189458 57634
rect 186313 57624 189458 57626
rect 186313 57568 186318 57624
rect 186374 57568 189458 57624
rect 186313 57566 189458 57568
rect 437473 57626 437539 57629
rect 437473 57624 440066 57626
rect 437473 57568 437478 57624
rect 437534 57568 440066 57624
rect 437473 57566 440066 57568
rect 186313 57563 186379 57566
rect 437473 57563 437539 57566
rect 440006 57324 440066 57566
rect 132217 57218 132283 57221
rect 130518 57216 132283 57218
rect 130518 57190 132222 57216
rect 129904 57160 132222 57190
rect 132278 57160 132283 57216
rect 129904 57158 132283 57160
rect 129904 57130 130578 57158
rect 132217 57155 132283 57158
rect 131205 56674 131271 56677
rect 130518 56672 131271 56674
rect 130518 56646 131210 56672
rect 129904 56616 131210 56646
rect 131266 56616 131271 56672
rect 129904 56614 131271 56616
rect 129904 56586 130578 56614
rect 131205 56611 131271 56614
rect 412173 56538 412239 56541
rect 409860 56536 412239 56538
rect 409860 56480 412178 56536
rect 412234 56480 412239 56536
rect 409860 56478 412239 56480
rect 412173 56475 412239 56478
rect 189398 56410 190072 56470
rect 187233 56402 187299 56405
rect 189398 56402 189458 56410
rect 187233 56400 189458 56402
rect 187233 56344 187238 56400
rect 187294 56344 189458 56400
rect 187233 56342 189458 56344
rect 187233 56339 187299 56342
rect 131205 56130 131271 56133
rect 130518 56128 131271 56130
rect 130518 56102 131210 56128
rect 129904 56072 131210 56102
rect 131266 56072 131271 56128
rect 129904 56070 131271 56072
rect 129904 56042 130578 56070
rect 131205 56067 131271 56070
rect 437473 56130 437539 56133
rect 437473 56128 440066 56130
rect 437473 56072 437478 56128
rect 437534 56072 440066 56128
rect 437473 56070 440066 56072
rect 437473 56067 437539 56070
rect 440006 55692 440066 56070
rect 131113 55450 131179 55453
rect 130518 55448 131179 55450
rect 130518 55422 131118 55448
rect 129904 55392 131118 55422
rect 131174 55392 131179 55448
rect 129904 55390 131179 55392
rect 129904 55362 130578 55390
rect 131113 55387 131179 55390
rect 189398 55322 190072 55382
rect 186313 55314 186379 55317
rect 189398 55314 189458 55322
rect 186313 55312 189458 55314
rect 186313 55256 186318 55312
rect 186374 55256 189458 55312
rect 186313 55254 189458 55256
rect 186313 55251 186379 55254
rect 132125 54906 132191 54909
rect 130518 54904 132191 54906
rect 130518 54878 132130 54904
rect 129904 54848 132130 54878
rect 132186 54848 132191 54904
rect 129904 54846 132191 54848
rect 129904 54818 130578 54846
rect 132125 54843 132191 54846
rect 411253 54634 411319 54637
rect 409860 54632 411319 54634
rect 409860 54576 411258 54632
rect 411314 54576 411319 54632
rect 409860 54574 411319 54576
rect 411253 54571 411319 54574
rect 437749 54634 437815 54637
rect 437749 54632 440066 54634
rect 437749 54576 437754 54632
rect 437810 54576 440066 54632
rect 437749 54574 440066 54576
rect 437749 54571 437815 54574
rect 131205 54362 131271 54365
rect 130518 54360 131271 54362
rect 130518 54334 131210 54360
rect 129904 54304 131210 54334
rect 131266 54304 131271 54360
rect 129904 54302 131271 54304
rect 129904 54274 130578 54302
rect 131205 54299 131271 54302
rect 189398 54234 190072 54294
rect 186313 54226 186379 54229
rect 189398 54226 189458 54234
rect 186313 54224 189458 54226
rect 186313 54168 186318 54224
rect 186374 54168 189458 54224
rect 440006 54196 440066 54574
rect 186313 54166 189458 54168
rect 186313 54163 186379 54166
rect 131205 53682 131271 53685
rect 130518 53680 131271 53682
rect 130518 53654 131210 53680
rect 129904 53624 131210 53654
rect 131266 53624 131271 53680
rect 129904 53622 131271 53624
rect 129904 53594 130578 53622
rect 131205 53619 131271 53622
rect 131665 53138 131731 53141
rect 130518 53136 131731 53138
rect 130518 53110 131670 53136
rect 129904 53080 131670 53110
rect 131726 53080 131731 53136
rect 129904 53078 131731 53080
rect 129904 53050 130578 53078
rect 131665 53075 131731 53078
rect 437473 53138 437539 53141
rect 437473 53136 440066 53138
rect 437473 53080 437478 53136
rect 437534 53080 440066 53136
rect 437473 53078 440066 53080
rect 437473 53075 437539 53078
rect 189398 53010 190072 53070
rect 187325 53002 187391 53005
rect 189398 53002 189458 53010
rect 187325 53000 189458 53002
rect 187325 52944 187330 53000
rect 187386 52944 189458 53000
rect 187325 52942 189458 52944
rect 187325 52939 187391 52942
rect 131113 52594 131179 52597
rect 411253 52594 411319 52597
rect 130518 52592 131179 52594
rect 130518 52566 131118 52592
rect 129904 52536 131118 52566
rect 131174 52536 131179 52592
rect 129904 52534 131179 52536
rect 409860 52592 411319 52594
rect 409860 52536 411258 52592
rect 411314 52536 411319 52592
rect 440006 52564 440066 53078
rect 543181 52730 543247 52733
rect 539948 52728 543247 52730
rect 539948 52672 543186 52728
rect 543242 52672 543247 52728
rect 539948 52670 543247 52672
rect 543181 52667 543247 52670
rect 409860 52534 411319 52536
rect 129904 52506 130578 52534
rect 131113 52531 131179 52534
rect 411253 52531 411319 52534
rect 132217 52050 132283 52053
rect 130518 52048 132283 52050
rect 130518 52022 132222 52048
rect 129904 51992 132222 52022
rect 132278 51992 132283 52048
rect 129904 51990 132283 51992
rect 129904 51962 130578 51990
rect 132217 51987 132283 51990
rect 189398 51922 190072 51982
rect 186313 51914 186379 51917
rect 189398 51914 189458 51922
rect 186313 51912 189458 51914
rect 186313 51856 186318 51912
rect 186374 51856 189458 51912
rect 186313 51854 189458 51856
rect 186313 51851 186379 51854
rect 437473 51642 437539 51645
rect 437473 51640 440066 51642
rect 437473 51584 437478 51640
rect 437534 51584 440066 51640
rect 437473 51582 440066 51584
rect 437473 51579 437539 51582
rect 131205 51370 131271 51373
rect 130518 51368 131271 51370
rect 130518 51342 131210 51368
rect 129904 51312 131210 51342
rect 131266 51312 131271 51368
rect 129904 51310 131271 51312
rect 129904 51282 130578 51310
rect 131205 51307 131271 51310
rect 440006 51068 440066 51582
rect 189398 50834 190072 50894
rect 132125 50826 132191 50829
rect 130518 50824 132191 50826
rect 130518 50798 132130 50824
rect 129904 50768 132130 50798
rect 132186 50768 132191 50824
rect 129904 50766 132191 50768
rect 129904 50738 130578 50766
rect 132125 50763 132191 50766
rect 186313 50826 186379 50829
rect 189398 50826 189458 50834
rect 186313 50824 189458 50826
rect 186313 50768 186318 50824
rect 186374 50768 189458 50824
rect 186313 50766 189458 50768
rect 186313 50763 186379 50766
rect 412449 50690 412515 50693
rect 409860 50688 412515 50690
rect 409860 50632 412454 50688
rect 412510 50632 412515 50688
rect 409860 50630 412515 50632
rect 412449 50627 412515 50630
rect 131849 50282 131915 50285
rect 130518 50280 131915 50282
rect 130518 50254 131854 50280
rect 129904 50224 131854 50254
rect 131910 50224 131915 50280
rect 129904 50222 131915 50224
rect 129904 50194 130578 50222
rect 131849 50219 131915 50222
rect 189398 49746 190072 49806
rect 186957 49738 187023 49741
rect 189398 49738 189458 49746
rect 186957 49736 189458 49738
rect 186957 49680 186962 49736
rect 187018 49680 189458 49736
rect 186957 49678 189458 49680
rect 186957 49675 187023 49678
rect 131205 49602 131271 49605
rect 130518 49600 131271 49602
rect 130518 49574 131210 49600
rect 129904 49544 131210 49574
rect 131266 49544 131271 49600
rect 129904 49542 131271 49544
rect 129904 49514 130578 49542
rect 131205 49539 131271 49542
rect 436829 49602 436895 49605
rect 436829 49600 440066 49602
rect 436829 49544 436834 49600
rect 436890 49544 440066 49600
rect 436829 49542 440066 49544
rect 436829 49539 436895 49542
rect 440006 49436 440066 49542
rect 131297 49058 131363 49061
rect 130518 49056 131363 49058
rect 130518 49030 131302 49056
rect 129904 49000 131302 49030
rect 131358 49000 131363 49056
rect 129904 48998 131363 49000
rect 129904 48970 130578 48998
rect 131297 48995 131363 48998
rect 411253 48786 411319 48789
rect 409860 48784 411319 48786
rect 409860 48728 411258 48784
rect 411314 48728 411319 48784
rect 409860 48726 411319 48728
rect 411253 48723 411319 48726
rect 189398 48522 190072 48582
rect 132309 48514 132375 48517
rect 130518 48512 132375 48514
rect 130518 48486 132314 48512
rect 129904 48456 132314 48486
rect 132370 48456 132375 48512
rect 129904 48454 132375 48456
rect 129904 48426 130578 48454
rect 132309 48451 132375 48454
rect 186313 48514 186379 48517
rect 189398 48514 189458 48522
rect 186313 48512 189458 48514
rect 186313 48456 186318 48512
rect 186374 48456 189458 48512
rect 186313 48454 189458 48456
rect 186313 48451 186379 48454
rect 437473 48242 437539 48245
rect 437473 48240 440066 48242
rect 437473 48184 437478 48240
rect 437534 48184 440066 48240
rect 437473 48182 440066 48184
rect 437473 48179 437539 48182
rect 440006 47940 440066 48182
rect 132217 47834 132283 47837
rect 130518 47832 132283 47834
rect 130518 47806 132222 47832
rect 129904 47776 132222 47806
rect 132278 47776 132283 47832
rect 129904 47774 132283 47776
rect 129904 47746 130578 47774
rect 132217 47771 132283 47774
rect 189398 47434 190072 47494
rect 186313 47426 186379 47429
rect 189398 47426 189458 47434
rect 186313 47424 189458 47426
rect 186313 47368 186318 47424
rect 186374 47368 189458 47424
rect 186313 47366 189458 47368
rect 186313 47363 186379 47366
rect 131205 47290 131271 47293
rect 130518 47288 131271 47290
rect 130518 47262 131210 47288
rect 129904 47232 131210 47262
rect 131266 47232 131271 47288
rect 129904 47230 131271 47232
rect 129904 47202 130578 47230
rect 131205 47227 131271 47230
rect 132401 46746 132467 46749
rect 412541 46746 412607 46749
rect 130518 46744 132467 46746
rect 130518 46718 132406 46744
rect 129904 46688 132406 46718
rect 132462 46688 132467 46744
rect 129904 46686 132467 46688
rect 409860 46744 412607 46746
rect 409860 46688 412546 46744
rect 412602 46688 412607 46744
rect 409860 46686 412607 46688
rect 129904 46658 130578 46686
rect 132401 46683 132467 46686
rect 412541 46683 412607 46686
rect 437473 46610 437539 46613
rect 437473 46608 440066 46610
rect 437473 46552 437478 46608
rect 437534 46552 440066 46608
rect 437473 46550 440066 46552
rect 437473 46547 437539 46550
rect 189398 46346 190072 46406
rect 187141 46338 187207 46341
rect 189398 46338 189458 46346
rect 187141 46336 189458 46338
rect 187141 46280 187146 46336
rect 187202 46280 189458 46336
rect 440006 46308 440066 46550
rect 580533 46338 580599 46341
rect 583520 46338 584960 46428
rect 580533 46336 584960 46338
rect 187141 46278 189458 46280
rect 580533 46280 580538 46336
rect 580594 46280 584960 46336
rect 580533 46278 584960 46280
rect 187141 46275 187207 46278
rect 580533 46275 580599 46278
rect 131113 46202 131179 46205
rect 130518 46200 131179 46202
rect 130518 46174 131118 46200
rect 129904 46144 131118 46174
rect 131174 46144 131179 46200
rect 583520 46188 584960 46278
rect 129904 46142 131179 46144
rect 129904 46114 130578 46142
rect 131113 46139 131179 46142
rect -960 45372 480 45612
rect 131205 45522 131271 45525
rect 130518 45520 131271 45522
rect 130518 45494 131210 45520
rect 129904 45464 131210 45494
rect 131266 45464 131271 45520
rect 129904 45462 131271 45464
rect 129904 45434 130578 45462
rect 131205 45459 131271 45462
rect 437473 45250 437539 45253
rect 437473 45248 440066 45250
rect 437473 45192 437478 45248
rect 437534 45192 440066 45248
rect 437473 45190 440066 45192
rect 437473 45187 437539 45190
rect 189398 45122 190072 45182
rect 186589 45114 186655 45117
rect 189398 45114 189458 45122
rect 186589 45112 189458 45114
rect 186589 45056 186594 45112
rect 186650 45056 189458 45112
rect 186589 45054 189458 45056
rect 186589 45051 186655 45054
rect 131941 44978 132007 44981
rect 130518 44976 132007 44978
rect 130518 44950 131946 44976
rect 129904 44920 131946 44950
rect 132002 44920 132007 44976
rect 129904 44918 132007 44920
rect 129904 44890 130578 44918
rect 131941 44915 132007 44918
rect 412265 44842 412331 44845
rect 409860 44840 412331 44842
rect 409860 44784 412270 44840
rect 412326 44784 412331 44840
rect 440006 44812 440066 45190
rect 409860 44782 412331 44784
rect 412265 44779 412331 44782
rect 131113 44434 131179 44437
rect 130518 44432 131179 44434
rect 130518 44406 131118 44432
rect 129904 44376 131118 44406
rect 131174 44376 131179 44432
rect 129904 44374 131179 44376
rect 129904 44346 130578 44374
rect 131113 44371 131179 44374
rect 189398 44034 190072 44094
rect 186405 44026 186471 44029
rect 189398 44026 189458 44034
rect 186405 44024 189458 44026
rect 186405 43968 186410 44024
rect 186466 43968 189458 44024
rect 186405 43966 189458 43968
rect 186405 43963 186471 43966
rect 131205 43754 131271 43757
rect 130518 43752 131271 43754
rect 130518 43726 131210 43752
rect 129904 43696 131210 43726
rect 131266 43696 131271 43752
rect 129904 43694 131271 43696
rect 129904 43666 130578 43694
rect 131205 43691 131271 43694
rect 437473 43618 437539 43621
rect 542997 43618 543063 43621
rect 437473 43616 440066 43618
rect 437473 43560 437478 43616
rect 437534 43560 440066 43616
rect 437473 43558 440066 43560
rect 539948 43616 543063 43618
rect 539948 43560 543002 43616
rect 543058 43560 543063 43616
rect 539948 43558 543063 43560
rect 437473 43555 437539 43558
rect 132033 43210 132099 43213
rect 130518 43208 132099 43210
rect 130518 43182 132038 43208
rect 129904 43152 132038 43182
rect 132094 43152 132099 43208
rect 440006 43180 440066 43558
rect 542997 43555 543063 43558
rect 129904 43150 132099 43152
rect 129904 43122 130578 43150
rect 132033 43147 132099 43150
rect 189398 42946 190072 43006
rect 186313 42938 186379 42941
rect 189398 42938 189458 42946
rect 186313 42936 189458 42938
rect 186313 42880 186318 42936
rect 186374 42880 189458 42936
rect 186313 42878 189458 42880
rect 186313 42875 186379 42878
rect 411253 42802 411319 42805
rect 409860 42800 411319 42802
rect 409860 42744 411258 42800
rect 411314 42744 411319 42800
rect 409860 42742 411319 42744
rect 411253 42739 411319 42742
rect 131205 42666 131271 42669
rect 130518 42664 131271 42666
rect 130518 42638 131210 42664
rect 129904 42608 131210 42638
rect 131266 42608 131271 42664
rect 129904 42606 131271 42608
rect 129904 42578 130578 42606
rect 131205 42603 131271 42606
rect 437473 42258 437539 42261
rect 437473 42256 440066 42258
rect 437473 42200 437478 42256
rect 437534 42200 440066 42256
rect 437473 42198 440066 42200
rect 437473 42195 437539 42198
rect 131113 41986 131179 41989
rect 130518 41984 131179 41986
rect 130518 41958 131118 41984
rect 129904 41928 131118 41958
rect 131174 41928 131179 41984
rect 129904 41926 131179 41928
rect 129904 41898 130578 41926
rect 131113 41923 131179 41926
rect 189398 41722 190072 41782
rect 186497 41714 186563 41717
rect 189398 41714 189458 41722
rect 186497 41712 189458 41714
rect 186497 41656 186502 41712
rect 186558 41656 189458 41712
rect 440006 41684 440066 42198
rect 186497 41654 189458 41656
rect 186497 41651 186563 41654
rect 132125 41442 132191 41445
rect 130150 41440 132191 41442
rect 130150 41408 132130 41440
rect 129904 41384 132130 41408
rect 132186 41384 132191 41440
rect 129904 41382 132191 41384
rect 129904 41348 130210 41382
rect 132125 41379 132191 41382
rect 131205 40898 131271 40901
rect 411253 40898 411319 40901
rect 130518 40896 131271 40898
rect 130518 40870 131210 40896
rect 129904 40840 131210 40870
rect 131266 40840 131271 40896
rect 129904 40838 131271 40840
rect 409860 40896 411319 40898
rect 409860 40840 411258 40896
rect 411314 40840 411319 40896
rect 409860 40838 411319 40840
rect 129904 40810 130578 40838
rect 131205 40835 131271 40838
rect 411253 40835 411319 40838
rect 189398 40634 190072 40694
rect 187233 40626 187299 40629
rect 189398 40626 189458 40634
rect 187233 40624 189458 40626
rect 187233 40568 187238 40624
rect 187294 40568 189458 40624
rect 187233 40566 189458 40568
rect 437473 40626 437539 40629
rect 437473 40624 440066 40626
rect 437473 40568 437478 40624
rect 437534 40568 440066 40624
rect 437473 40566 440066 40568
rect 187233 40563 187299 40566
rect 437473 40563 437539 40566
rect 131113 40354 131179 40357
rect 130518 40352 131179 40354
rect 130518 40326 131118 40352
rect 129904 40296 131118 40326
rect 131174 40296 131179 40352
rect 129904 40294 131179 40296
rect 129904 40266 130578 40294
rect 131113 40291 131179 40294
rect 440006 40052 440066 40566
rect 131849 39674 131915 39677
rect 130518 39672 131915 39674
rect 130518 39646 131854 39672
rect 129904 39616 131854 39646
rect 131910 39616 131915 39672
rect 129904 39614 131915 39616
rect 129904 39586 130578 39614
rect 131849 39611 131915 39614
rect 189398 39546 190072 39606
rect 186957 39538 187023 39541
rect 189398 39538 189458 39546
rect 186957 39536 189458 39538
rect 186957 39480 186962 39536
rect 187018 39480 189458 39536
rect 186957 39478 189458 39480
rect 186957 39475 187023 39478
rect 132493 39130 132559 39133
rect 130518 39128 132559 39130
rect 130518 39102 132498 39128
rect 129904 39072 132498 39102
rect 132554 39072 132559 39128
rect 129904 39070 132559 39072
rect 129904 39042 130578 39070
rect 132493 39067 132559 39070
rect 411253 38858 411319 38861
rect 409860 38856 411319 38858
rect 409860 38800 411258 38856
rect 411314 38800 411319 38856
rect 409860 38798 411319 38800
rect 411253 38795 411319 38798
rect 131205 38586 131271 38589
rect 130518 38584 131271 38586
rect 130518 38558 131210 38584
rect 129904 38528 131210 38558
rect 131266 38528 131271 38584
rect 129904 38526 131271 38528
rect 129904 38498 130578 38526
rect 131205 38523 131271 38526
rect 189398 38458 190072 38518
rect 186405 38450 186471 38453
rect 189398 38450 189458 38458
rect 186405 38448 189458 38450
rect 186405 38392 186410 38448
rect 186466 38392 189458 38448
rect 186405 38390 189458 38392
rect 437473 38450 437539 38453
rect 440006 38450 440066 38556
rect 437473 38448 440066 38450
rect 437473 38392 437478 38448
rect 437534 38392 440066 38448
rect 437473 38390 440066 38392
rect 186405 38387 186471 38390
rect 437473 38387 437539 38390
rect 131113 37906 131179 37909
rect 130518 37904 131179 37906
rect 130518 37878 131118 37904
rect 129904 37848 131118 37878
rect 131174 37848 131179 37904
rect 129904 37846 131179 37848
rect 129904 37818 130578 37846
rect 131113 37843 131179 37846
rect 131665 37362 131731 37365
rect 130518 37360 131731 37362
rect 130518 37334 131670 37360
rect 129904 37304 131670 37334
rect 131726 37304 131731 37360
rect 129904 37302 131731 37304
rect 129904 37274 130578 37302
rect 131665 37299 131731 37302
rect 186313 37362 186379 37365
rect 186313 37360 189642 37362
rect 186313 37304 186318 37360
rect 186374 37334 189642 37360
rect 186374 37304 190164 37334
rect 186313 37302 190164 37304
rect 186313 37299 186379 37302
rect 189582 37274 190164 37302
rect 437473 37226 437539 37229
rect 437473 37224 440066 37226
rect 437473 37168 437478 37224
rect 437534 37168 440066 37224
rect 437473 37166 440066 37168
rect 437473 37163 437539 37166
rect 411253 36954 411319 36957
rect 409860 36952 411319 36954
rect 409860 36896 411258 36952
rect 411314 36896 411319 36952
rect 440006 36924 440066 37166
rect 409860 36894 411319 36896
rect 411253 36891 411319 36894
rect 131297 36818 131363 36821
rect 130518 36816 131363 36818
rect 130518 36790 131302 36816
rect 129904 36760 131302 36790
rect 131358 36760 131363 36816
rect 129904 36758 131363 36760
rect 129904 36730 130578 36758
rect 131297 36755 131363 36758
rect 189398 36146 190072 36206
rect 131205 36138 131271 36141
rect 130518 36136 131271 36138
rect 130518 36110 131210 36136
rect 129904 36080 131210 36110
rect 131266 36080 131271 36136
rect 129904 36078 131271 36080
rect 129904 36050 130578 36078
rect 131205 36075 131271 36078
rect 186313 36138 186379 36141
rect 189398 36138 189458 36146
rect 186313 36136 189458 36138
rect 186313 36080 186318 36136
rect 186374 36080 189458 36136
rect 186313 36078 189458 36080
rect 186313 36075 186379 36078
rect 437473 35866 437539 35869
rect 437473 35864 440066 35866
rect 437473 35808 437478 35864
rect 437534 35808 440066 35864
rect 437473 35806 440066 35808
rect 437473 35803 437539 35806
rect 131205 35594 131271 35597
rect 130518 35592 131271 35594
rect 130518 35566 131210 35592
rect 129904 35536 131210 35566
rect 131266 35536 131271 35592
rect 129904 35534 131271 35536
rect 129904 35506 130578 35534
rect 131205 35531 131271 35534
rect 440006 35428 440066 35806
rect 189398 35058 190072 35118
rect 131113 35050 131179 35053
rect 130518 35048 131179 35050
rect 130518 35022 131118 35048
rect 129904 34992 131118 35022
rect 131174 34992 131179 35048
rect 129904 34990 131179 34992
rect 129904 34962 130578 34990
rect 131113 34987 131179 34990
rect 186405 35050 186471 35053
rect 189398 35050 189458 35058
rect 186405 35048 189458 35050
rect 186405 34992 186410 35048
rect 186466 34992 189458 35048
rect 186405 34990 189458 34992
rect 186405 34987 186471 34990
rect 411253 34914 411319 34917
rect 409860 34912 411319 34914
rect 409860 34856 411258 34912
rect 411314 34856 411319 34912
rect 409860 34854 411319 34856
rect 411253 34851 411319 34854
rect 543089 34642 543155 34645
rect 539948 34640 543155 34642
rect 539948 34584 543094 34640
rect 543150 34584 543155 34640
rect 539948 34582 543155 34584
rect 543089 34579 543155 34582
rect 132125 34506 132191 34509
rect 130518 34504 132191 34506
rect 130518 34478 132130 34504
rect 129904 34448 132130 34478
rect 132186 34448 132191 34504
rect 129904 34446 132191 34448
rect 129904 34418 130578 34446
rect 132125 34443 132191 34446
rect 437473 34098 437539 34101
rect 437473 34096 440066 34098
rect 437473 34040 437478 34096
rect 437534 34040 440066 34096
rect 437473 34038 440066 34040
rect 437473 34035 437539 34038
rect 189398 33834 190072 33894
rect 132033 33826 132099 33829
rect 130518 33824 132099 33826
rect 130518 33798 132038 33824
rect 129904 33768 132038 33798
rect 132094 33768 132099 33824
rect 129904 33766 132099 33768
rect 129904 33738 130578 33766
rect 132033 33763 132099 33766
rect 186313 33826 186379 33829
rect 189398 33826 189458 33834
rect 186313 33824 189458 33826
rect 186313 33768 186318 33824
rect 186374 33768 189458 33824
rect 440006 33796 440066 34038
rect 186313 33766 189458 33768
rect 186313 33763 186379 33766
rect 132217 33282 132283 33285
rect 130518 33280 132283 33282
rect 130518 33254 132222 33280
rect 129904 33224 132222 33254
rect 132278 33224 132283 33280
rect 129904 33222 132283 33224
rect 129904 33194 130578 33222
rect 132217 33219 132283 33222
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 411253 33010 411319 33013
rect 409860 33008 411319 33010
rect 409860 32952 411258 33008
rect 411314 32952 411319 33008
rect 583520 32996 584960 33086
rect 409860 32950 411319 32952
rect 411253 32947 411319 32950
rect 189398 32746 190072 32806
rect 131205 32738 131271 32741
rect 130518 32736 131271 32738
rect 130518 32710 131210 32736
rect 129904 32680 131210 32710
rect 131266 32680 131271 32736
rect 129904 32678 131271 32680
rect 129904 32650 130578 32678
rect 131205 32675 131271 32678
rect 186405 32738 186471 32741
rect 189398 32738 189458 32746
rect 186405 32736 189458 32738
rect 186405 32680 186410 32736
rect 186466 32680 189458 32736
rect 186405 32678 189458 32680
rect 437473 32738 437539 32741
rect 437473 32736 440066 32738
rect 437473 32680 437478 32736
rect 437534 32680 440066 32736
rect 437473 32678 440066 32680
rect 186405 32675 186471 32678
rect 437473 32675 437539 32678
rect -960 32316 480 32556
rect 440006 32300 440066 32678
rect 131113 32058 131179 32061
rect 130518 32056 131179 32058
rect 130518 32030 131118 32056
rect 129904 32000 131118 32030
rect 131174 32000 131179 32056
rect 129904 31998 131179 32000
rect 129904 31970 130578 31998
rect 131113 31995 131179 31998
rect 186313 31786 186379 31789
rect 186313 31784 189826 31786
rect 186313 31728 186318 31784
rect 186374 31758 189826 31784
rect 186374 31728 190010 31758
rect 186313 31726 190010 31728
rect 186313 31723 186379 31726
rect 189766 31718 190010 31726
rect 189766 31698 190072 31718
rect 189950 31658 190072 31698
rect 131205 31514 131271 31517
rect 130518 31512 131271 31514
rect 130518 31486 131210 31512
rect 129904 31456 131210 31486
rect 131266 31456 131271 31512
rect 129904 31454 131271 31456
rect 129904 31426 130578 31454
rect 131205 31451 131271 31454
rect 437473 31242 437539 31245
rect 437473 31240 440066 31242
rect 437473 31184 437478 31240
rect 437534 31184 440066 31240
rect 437473 31182 440066 31184
rect 437473 31179 437539 31182
rect 411253 31106 411319 31109
rect 409860 31104 411319 31106
rect 409860 31048 411258 31104
rect 411314 31048 411319 31104
rect 409860 31046 411319 31048
rect 411253 31043 411319 31046
rect 131297 30970 131363 30973
rect 130518 30968 131363 30970
rect 130518 30942 131302 30968
rect 129904 30912 131302 30942
rect 131358 30912 131363 30968
rect 129904 30910 131363 30912
rect 129904 30882 130578 30910
rect 131297 30907 131363 30910
rect 440006 30804 440066 31182
rect 186313 30562 186379 30565
rect 190134 30562 190194 30668
rect 186313 30560 190194 30562
rect 186313 30504 186318 30560
rect 186374 30504 190194 30560
rect 186313 30502 190194 30504
rect 186313 30499 186379 30502
rect 131113 30426 131179 30429
rect 130150 30424 131179 30426
rect 129782 30290 129842 30396
rect 130150 30368 131118 30424
rect 131174 30368 131179 30424
rect 130150 30366 131179 30368
rect 130150 30290 130210 30366
rect 131113 30363 131179 30366
rect 129782 30230 130210 30290
rect 133137 28930 133203 28933
rect 405733 28930 405799 28933
rect 133137 28928 405799 28930
rect 133137 28872 133142 28928
rect 133198 28872 405738 28928
rect 405794 28872 405799 28928
rect 133137 28870 405799 28872
rect 133137 28867 133203 28870
rect 405733 28867 405799 28870
rect 131757 28794 131823 28797
rect 397453 28794 397519 28797
rect 131757 28792 397519 28794
rect 131757 28736 131762 28792
rect 131818 28736 397458 28792
rect 397514 28736 397519 28792
rect 131757 28734 397519 28736
rect 131757 28731 131823 28734
rect 397453 28731 397519 28734
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19260 480 19500
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6340 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 583520 6476 584960 6566
<< via3 >>
rect 239654 299780 239718 299844
rect 243054 299704 243118 299708
rect 243054 299648 243082 299704
rect 243082 299648 243118 299704
rect 243054 299644 243118 299648
rect 55854 299568 55918 299572
rect 55854 299512 55862 299568
rect 55862 299512 55918 299568
rect 55854 299508 55918 299512
rect 73660 298148 73724 298212
rect 77892 298148 77956 298212
rect 81756 298148 81820 298212
rect 85436 298148 85500 298212
rect 91876 298148 91940 298212
rect 95556 298148 95620 298212
rect 95924 298148 95988 298212
rect 99420 298148 99484 298212
rect 102916 298148 102980 298212
rect 103284 298208 103348 298212
rect 103284 298152 103298 298208
rect 103298 298152 103348 298208
rect 103284 298148 103348 298152
rect 225460 298148 225524 298212
rect 229140 298148 229204 298212
rect 257844 298148 257908 298212
rect 65564 298012 65628 298076
rect 66668 298012 66732 298076
rect 67772 298072 67836 298076
rect 67772 298016 67822 298072
rect 67822 298016 67836 298072
rect 67772 298012 67836 298016
rect 69244 298012 69308 298076
rect 70164 298072 70228 298076
rect 70164 298016 70214 298072
rect 70214 298016 70228 298072
rect 70164 298012 70228 298016
rect 71452 298072 71516 298076
rect 71452 298016 71502 298072
rect 71502 298016 71516 298072
rect 71452 298012 71516 298016
rect 72556 298012 72620 298076
rect 75132 298012 75196 298076
rect 76236 298012 76300 298076
rect 77156 298072 77220 298076
rect 77156 298016 77170 298072
rect 77170 298016 77220 298072
rect 77156 298012 77220 298016
rect 78260 298012 78324 298076
rect 79364 298012 79428 298076
rect 80836 298012 80900 298076
rect 82124 298012 82188 298076
rect 83228 298012 83292 298076
rect 84516 298012 84580 298076
rect 86540 298012 86604 298076
rect 87828 298012 87892 298076
rect 89300 298012 89364 298076
rect 90772 298012 90836 298076
rect 93164 298012 93228 298076
rect 93532 298012 93596 298076
rect 94452 298012 94516 298076
rect 79732 297936 79796 297940
rect 79732 297880 79782 297936
rect 79782 297880 79796 297936
rect 79732 297876 79796 297880
rect 80284 297876 80348 297940
rect 83044 297876 83108 297940
rect 86908 297876 86972 297940
rect 87644 297876 87708 297940
rect 88932 297876 88996 297940
rect 90220 297876 90284 297940
rect 91324 297876 91388 297940
rect 92612 297876 92676 297940
rect 95004 297876 95068 297940
rect 96660 298072 96724 298076
rect 96660 298016 96710 298072
rect 96710 298016 96724 298072
rect 96660 298012 96724 298016
rect 97948 298012 98012 298076
rect 99052 298012 99116 298076
rect 97028 297876 97092 297940
rect 98316 297876 98380 297940
rect 100524 298072 100588 298076
rect 100524 298016 100574 298072
rect 100574 298016 100588 298072
rect 100524 298012 100588 298016
rect 101812 298072 101876 298076
rect 101812 298016 101862 298072
rect 101862 298016 101876 298072
rect 101812 298012 101876 298016
rect 104388 298012 104452 298076
rect 105676 298012 105740 298076
rect 106596 298012 106660 298076
rect 106964 298012 107028 298076
rect 107884 298012 107948 298076
rect 109356 298012 109420 298076
rect 110644 298012 110708 298076
rect 113036 298072 113100 298076
rect 113036 298016 113050 298072
rect 113050 298016 113100 298072
rect 113036 298012 113100 298016
rect 114324 298012 114388 298076
rect 115612 298012 115676 298076
rect 116900 298012 116964 298076
rect 215892 298072 215956 298076
rect 261524 298148 261588 298212
rect 261892 298148 261956 298212
rect 265204 298148 265268 298212
rect 271828 298148 271892 298212
rect 275508 298148 275572 298212
rect 215892 298016 215906 298072
rect 215906 298016 215956 298072
rect 215892 298012 215956 298016
rect 226748 298012 226812 298076
rect 227852 298012 227916 298076
rect 231348 298012 231412 298076
rect 232636 298012 232700 298076
rect 233556 298012 233620 298076
rect 235028 298012 235092 298076
rect 237236 298072 237300 298076
rect 237236 298016 237250 298072
rect 237250 298016 237300 298072
rect 237236 298012 237300 298016
rect 239260 298012 239324 298076
rect 240364 298012 240428 298076
rect 240732 298012 240796 298076
rect 242940 298072 243004 298076
rect 242940 298016 242954 298072
rect 242954 298016 243004 298072
rect 242940 298012 243004 298016
rect 244044 298072 244108 298076
rect 244044 298016 244094 298072
rect 244094 298016 244108 298072
rect 244044 298012 244108 298016
rect 244412 298012 244476 298076
rect 245516 298072 245580 298076
rect 245516 298016 245566 298072
rect 245566 298016 245580 298072
rect 245516 298012 245580 298016
rect 246804 298072 246868 298076
rect 246804 298016 246854 298072
rect 246854 298016 246868 298072
rect 246804 298012 246868 298016
rect 247908 298012 247972 298076
rect 249380 298012 249444 298076
rect 250668 298012 250732 298076
rect 252508 298012 252572 298076
rect 253612 298012 253676 298076
rect 254900 298012 254964 298076
rect 256004 298012 256068 298076
rect 257108 298012 257172 298076
rect 259316 298012 259380 298076
rect 260788 298012 260852 298076
rect 101444 297876 101508 297940
rect 104020 297876 104084 297940
rect 105308 297876 105372 297940
rect 107700 297876 107764 297940
rect 111932 297876 111996 297940
rect 237788 297876 237852 297940
rect 242020 297876 242084 297940
rect 246620 297876 246684 297940
rect 247724 297876 247788 297940
rect 249012 297876 249076 297940
rect 250300 297876 250364 297940
rect 251404 297876 251468 297940
rect 253060 297876 253124 297940
rect 254532 297876 254596 297940
rect 255636 297876 255700 297940
rect 256740 297876 256804 297940
rect 259132 297876 259196 297940
rect 260604 297876 260668 297940
rect 263180 298012 263244 298076
rect 274404 298012 274468 298076
rect 276796 298012 276860 298076
rect 262996 297876 263060 297940
rect 85804 297740 85868 297804
rect 100708 297740 100772 297804
rect 236500 297740 236564 297804
rect 241836 297740 241900 297804
rect 245700 297740 245764 297804
rect 251956 297740 252020 297804
rect 258396 297740 258460 297804
rect 267964 297468 268028 297532
rect 230060 297196 230124 297260
rect 83964 297060 84028 297124
rect 266676 297060 266740 297124
rect 264100 296924 264164 296988
rect 266860 296924 266924 296988
rect 238340 296788 238404 296852
rect 264468 296788 264532 296852
rect 265756 296788 265820 296852
rect 267596 296788 267660 296852
rect 269252 296788 269316 296852
rect 270540 296788 270604 296852
rect 273116 296848 273180 296852
rect 273116 296792 273130 296848
rect 273130 296792 273180 296848
rect 273116 296788 273180 296792
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 132000 31574 140058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 132000 38414 146898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 132000 42134 150618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 381500 49574 410058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381500 56414 416898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 381500 60134 384618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 381500 63854 388338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 381500 67574 392058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 381500 74414 398898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 381500 78134 402618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 381500 81854 406338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 381500 85574 410058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381500 92414 416898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 381500 96134 384618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 381500 99854 388338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 381500 103574 392058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 381500 110414 398898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 381500 114134 402618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 381500 117854 406338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 381500 121574 410058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381500 128414 416898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 381500 132134 384618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 381500 135854 388338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 381500 139574 392058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 381500 146414 398898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 50952 363454 51300 363486
rect 50952 363218 51008 363454
rect 51244 363218 51300 363454
rect 50952 363134 51300 363218
rect 50952 362898 51008 363134
rect 51244 362898 51300 363134
rect 50952 362866 51300 362898
rect 144656 363454 145004 363486
rect 144656 363218 144712 363454
rect 144948 363218 145004 363454
rect 144656 363134 145004 363218
rect 144656 362898 144712 363134
rect 144948 362898 145004 363134
rect 144656 362866 145004 362898
rect 50272 345454 50620 345486
rect 50272 345218 50328 345454
rect 50564 345218 50620 345454
rect 50272 345134 50620 345218
rect 50272 344898 50328 345134
rect 50564 344898 50620 345134
rect 50272 344866 50620 344898
rect 145336 345454 145684 345486
rect 145336 345218 145392 345454
rect 145628 345218 145684 345454
rect 145336 345134 145684 345218
rect 145336 344898 145392 345134
rect 145628 344898 145684 345134
rect 145336 344866 145684 344898
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 50952 327454 51300 327486
rect 50952 327218 51008 327454
rect 51244 327218 51300 327454
rect 50952 327134 51300 327218
rect 50952 326898 51008 327134
rect 51244 326898 51300 327134
rect 50952 326866 51300 326898
rect 144656 327454 145004 327486
rect 144656 327218 144712 327454
rect 144948 327218 145004 327454
rect 144656 327134 145004 327218
rect 144656 326898 144712 327134
rect 144948 326898 145004 327134
rect 144656 326866 145004 326898
rect 50272 309454 50620 309486
rect 50272 309218 50328 309454
rect 50564 309218 50620 309454
rect 50272 309134 50620 309218
rect 50272 308898 50328 309134
rect 50564 308898 50620 309134
rect 50272 308866 50620 308898
rect 145336 309454 145684 309486
rect 145336 309218 145392 309454
rect 145628 309218 145684 309454
rect 145336 309134 145684 309218
rect 145336 308898 145392 309134
rect 145628 308898 145684 309134
rect 145336 308866 145684 308898
rect 55856 299573 55916 300106
rect 55853 299572 55919 299573
rect 55853 299508 55854 299572
rect 55918 299508 55919 299572
rect 65512 299570 65572 300106
rect 66736 299570 66796 300106
rect 67824 299570 67884 300106
rect 65512 299510 65626 299570
rect 55853 299507 55919 299508
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 65566 298077 65626 299510
rect 66670 299510 66796 299570
rect 67774 299510 67884 299570
rect 69184 299570 69244 300106
rect 70136 299570 70196 300106
rect 71360 299570 71420 300106
rect 72584 299570 72644 300106
rect 73672 299570 73732 300106
rect 69184 299510 69306 299570
rect 70136 299510 70226 299570
rect 71360 299510 71514 299570
rect 66670 298077 66730 299510
rect 67774 298077 67834 299510
rect 69246 298077 69306 299510
rect 70166 298077 70226 299510
rect 71454 298077 71514 299510
rect 72558 299510 72644 299570
rect 73662 299510 73732 299570
rect 75032 299570 75092 300106
rect 76120 299570 76180 300106
rect 77208 299570 77268 300106
rect 75032 299510 75194 299570
rect 76120 299510 76298 299570
rect 72558 298077 72618 299510
rect 73662 298213 73722 299510
rect 73659 298212 73725 298213
rect 73659 298148 73660 298212
rect 73724 298148 73725 298212
rect 73659 298147 73725 298148
rect 75134 298077 75194 299510
rect 76238 298077 76298 299510
rect 77158 299510 77268 299570
rect 77888 299570 77948 300106
rect 78296 299570 78356 300106
rect 77888 299510 77954 299570
rect 77158 298077 77218 299510
rect 77894 298213 77954 299510
rect 78262 299510 78356 299570
rect 79248 299570 79308 300106
rect 79656 299570 79716 300106
rect 80336 299570 80396 300106
rect 79248 299510 79426 299570
rect 79656 299510 79794 299570
rect 77891 298212 77957 298213
rect 77891 298148 77892 298212
rect 77956 298148 77957 298212
rect 77891 298147 77957 298148
rect 78262 298077 78322 299510
rect 79366 298077 79426 299510
rect 65563 298076 65629 298077
rect 65563 298012 65564 298076
rect 65628 298012 65629 298076
rect 65563 298011 65629 298012
rect 66667 298076 66733 298077
rect 66667 298012 66668 298076
rect 66732 298012 66733 298076
rect 66667 298011 66733 298012
rect 67771 298076 67837 298077
rect 67771 298012 67772 298076
rect 67836 298012 67837 298076
rect 67771 298011 67837 298012
rect 69243 298076 69309 298077
rect 69243 298012 69244 298076
rect 69308 298012 69309 298076
rect 69243 298011 69309 298012
rect 70163 298076 70229 298077
rect 70163 298012 70164 298076
rect 70228 298012 70229 298076
rect 70163 298011 70229 298012
rect 71451 298076 71517 298077
rect 71451 298012 71452 298076
rect 71516 298012 71517 298076
rect 71451 298011 71517 298012
rect 72555 298076 72621 298077
rect 72555 298012 72556 298076
rect 72620 298012 72621 298076
rect 72555 298011 72621 298012
rect 75131 298076 75197 298077
rect 75131 298012 75132 298076
rect 75196 298012 75197 298076
rect 75131 298011 75197 298012
rect 76235 298076 76301 298077
rect 76235 298012 76236 298076
rect 76300 298012 76301 298076
rect 76235 298011 76301 298012
rect 77155 298076 77221 298077
rect 77155 298012 77156 298076
rect 77220 298012 77221 298076
rect 77155 298011 77221 298012
rect 78259 298076 78325 298077
rect 78259 298012 78260 298076
rect 78324 298012 78325 298076
rect 78259 298011 78325 298012
rect 79363 298076 79429 298077
rect 79363 298012 79364 298076
rect 79428 298012 79429 298076
rect 79363 298011 79429 298012
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 132000 45854 154338
rect 48954 266614 49574 298000
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 132000 49574 158058
rect 55794 273454 56414 298000
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 132000 56414 164898
rect 59514 277174 60134 298000
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 132000 60134 132618
rect 63234 280894 63854 298000
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 132000 63854 136338
rect 66954 284614 67574 298000
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 132000 67574 140058
rect 73794 291454 74414 298000
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 132000 74414 146898
rect 77514 295174 78134 298000
rect 79734 297941 79794 299510
rect 80286 299510 80396 299570
rect 80744 299570 80804 300106
rect 81832 299570 81892 300106
rect 80744 299510 80898 299570
rect 80286 297941 80346 299510
rect 80838 298077 80898 299510
rect 81758 299510 81892 299570
rect 81968 299570 82028 300106
rect 83056 299570 83116 300106
rect 81968 299510 82186 299570
rect 81758 298213 81818 299510
rect 81755 298212 81821 298213
rect 81755 298148 81756 298212
rect 81820 298148 81821 298212
rect 81755 298147 81821 298148
rect 82126 298077 82186 299510
rect 83046 299510 83116 299570
rect 83192 299570 83252 300106
rect 84144 299570 84204 300106
rect 83192 299510 83290 299570
rect 80835 298076 80901 298077
rect 80835 298012 80836 298076
rect 80900 298012 80901 298076
rect 80835 298011 80901 298012
rect 82123 298076 82189 298077
rect 82123 298012 82124 298076
rect 82188 298012 82189 298076
rect 82123 298011 82189 298012
rect 79731 297940 79797 297941
rect 79731 297876 79732 297940
rect 79796 297876 79797 297940
rect 79731 297875 79797 297876
rect 80283 297940 80349 297941
rect 80283 297876 80284 297940
rect 80348 297876 80349 297940
rect 80283 297875 80349 297876
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 132000 78134 150618
rect 81234 262894 81854 298000
rect 83046 297941 83106 299510
rect 83230 298077 83290 299510
rect 83966 299510 84204 299570
rect 84416 299570 84476 300106
rect 85504 299570 85564 300106
rect 84416 299510 84578 299570
rect 83227 298076 83293 298077
rect 83227 298012 83228 298076
rect 83292 298012 83293 298076
rect 83227 298011 83293 298012
rect 83043 297940 83109 297941
rect 83043 297876 83044 297940
rect 83108 297876 83109 297940
rect 83043 297875 83109 297876
rect 83966 297125 84026 299510
rect 84518 298077 84578 299510
rect 85438 299510 85564 299570
rect 85640 299570 85700 300106
rect 86592 299570 86652 300106
rect 85640 299510 85866 299570
rect 85438 298213 85498 299510
rect 85435 298212 85501 298213
rect 85435 298148 85436 298212
rect 85500 298148 85501 298212
rect 85435 298147 85501 298148
rect 84515 298076 84581 298077
rect 84515 298012 84516 298076
rect 84580 298012 84581 298076
rect 84515 298011 84581 298012
rect 83963 297124 84029 297125
rect 83963 297060 83964 297124
rect 84028 297060 84029 297124
rect 83963 297059 84029 297060
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 132000 81854 154338
rect 84954 266614 85574 298000
rect 85806 297805 85866 299510
rect 86542 299510 86652 299570
rect 86864 299570 86924 300106
rect 87680 299570 87740 300106
rect 86864 299510 86970 299570
rect 86542 298077 86602 299510
rect 86539 298076 86605 298077
rect 86539 298012 86540 298076
rect 86604 298012 86605 298076
rect 86539 298011 86605 298012
rect 86910 297941 86970 299510
rect 87646 299510 87740 299570
rect 87816 299570 87876 300106
rect 88904 299570 88964 300106
rect 89312 299570 89372 300106
rect 90264 299570 90324 300106
rect 87816 299510 87890 299570
rect 88904 299510 88994 299570
rect 87646 297941 87706 299510
rect 87830 298077 87890 299510
rect 87827 298076 87893 298077
rect 87827 298012 87828 298076
rect 87892 298012 87893 298076
rect 87827 298011 87893 298012
rect 88934 297941 88994 299510
rect 89302 299510 89372 299570
rect 90222 299510 90324 299570
rect 90672 299570 90732 300106
rect 91352 299570 91412 300106
rect 91896 299570 91956 300106
rect 90672 299510 90834 299570
rect 89302 298077 89362 299510
rect 89299 298076 89365 298077
rect 89299 298012 89300 298076
rect 89364 298012 89365 298076
rect 89299 298011 89365 298012
rect 90222 297941 90282 299510
rect 90774 298077 90834 299510
rect 91326 299510 91412 299570
rect 91878 299510 91956 299570
rect 92440 299570 92500 300106
rect 93120 299570 93180 300106
rect 93528 299570 93588 300106
rect 94344 299842 94404 300106
rect 94888 299842 94948 300106
rect 94344 299782 94514 299842
rect 94888 299782 95066 299842
rect 92440 299510 92674 299570
rect 93120 299510 93226 299570
rect 93528 299510 93594 299570
rect 90771 298076 90837 298077
rect 90771 298012 90772 298076
rect 90836 298012 90837 298076
rect 90771 298011 90837 298012
rect 91326 297941 91386 299510
rect 91878 298213 91938 299510
rect 91875 298212 91941 298213
rect 91875 298148 91876 298212
rect 91940 298148 91941 298212
rect 91875 298147 91941 298148
rect 86907 297940 86973 297941
rect 86907 297876 86908 297940
rect 86972 297876 86973 297940
rect 86907 297875 86973 297876
rect 87643 297940 87709 297941
rect 87643 297876 87644 297940
rect 87708 297876 87709 297940
rect 87643 297875 87709 297876
rect 88931 297940 88997 297941
rect 88931 297876 88932 297940
rect 88996 297876 88997 297940
rect 88931 297875 88997 297876
rect 90219 297940 90285 297941
rect 90219 297876 90220 297940
rect 90284 297876 90285 297940
rect 90219 297875 90285 297876
rect 91323 297940 91389 297941
rect 91323 297876 91324 297940
rect 91388 297876 91389 297940
rect 91323 297875 91389 297876
rect 85803 297804 85869 297805
rect 85803 297740 85804 297804
rect 85868 297740 85869 297804
rect 85803 297739 85869 297740
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 132000 85574 158058
rect 91794 273454 92414 298000
rect 92614 297941 92674 299510
rect 93166 298077 93226 299510
rect 93534 298077 93594 299510
rect 94454 298077 94514 299782
rect 93163 298076 93229 298077
rect 93163 298012 93164 298076
rect 93228 298012 93229 298076
rect 93163 298011 93229 298012
rect 93531 298076 93597 298077
rect 93531 298012 93532 298076
rect 93596 298012 93597 298076
rect 93531 298011 93597 298012
rect 94451 298076 94517 298077
rect 94451 298012 94452 298076
rect 94516 298012 94517 298076
rect 94451 298011 94517 298012
rect 95006 297941 95066 299782
rect 95568 299570 95628 300106
rect 95976 299570 96036 300106
rect 95558 299510 95628 299570
rect 95926 299510 96036 299570
rect 96656 299570 96716 300106
rect 97064 299570 97124 300106
rect 97880 299842 97940 300106
rect 97880 299782 98010 299842
rect 96656 299510 96722 299570
rect 95558 298213 95618 299510
rect 95926 298213 95986 299510
rect 95555 298212 95621 298213
rect 95555 298148 95556 298212
rect 95620 298148 95621 298212
rect 95555 298147 95621 298148
rect 95923 298212 95989 298213
rect 95923 298148 95924 298212
rect 95988 298148 95989 298212
rect 95923 298147 95989 298148
rect 96662 298077 96722 299510
rect 97030 299510 97124 299570
rect 96659 298076 96725 298077
rect 96659 298012 96660 298076
rect 96724 298012 96725 298076
rect 96659 298011 96725 298012
rect 92611 297940 92677 297941
rect 92611 297876 92612 297940
rect 92676 297876 92677 297940
rect 92611 297875 92677 297876
rect 95003 297940 95069 297941
rect 95003 297876 95004 297940
rect 95068 297876 95069 297940
rect 95003 297875 95069 297876
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 132000 92414 164898
rect 95514 277174 96134 298000
rect 97030 297941 97090 299510
rect 97950 298077 98010 299782
rect 98288 299570 98348 300106
rect 99104 299570 99164 300106
rect 98288 299510 98378 299570
rect 97947 298076 98013 298077
rect 97947 298012 97948 298076
rect 98012 298012 98013 298076
rect 97947 298011 98013 298012
rect 98318 297941 98378 299510
rect 99054 299510 99164 299570
rect 99376 299570 99436 300106
rect 100600 299842 100660 300106
rect 100526 299782 100660 299842
rect 99376 299510 99482 299570
rect 99054 298077 99114 299510
rect 99422 298213 99482 299510
rect 99419 298212 99485 298213
rect 99419 298148 99420 298212
rect 99484 298148 99485 298212
rect 99419 298147 99485 298148
rect 100526 298077 100586 299782
rect 100736 299570 100796 300106
rect 100710 299510 100796 299570
rect 101416 299570 101476 300106
rect 101824 299570 101884 300106
rect 101416 299510 101506 299570
rect 99051 298076 99117 298077
rect 99051 298012 99052 298076
rect 99116 298012 99117 298076
rect 99051 298011 99117 298012
rect 100523 298076 100589 298077
rect 100523 298012 100524 298076
rect 100588 298012 100589 298076
rect 100523 298011 100589 298012
rect 97027 297940 97093 297941
rect 97027 297876 97028 297940
rect 97092 297876 97093 297940
rect 97027 297875 97093 297876
rect 98315 297940 98381 297941
rect 98315 297876 98316 297940
rect 98380 297876 98381 297940
rect 98315 297875 98381 297876
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 132000 96134 132618
rect 99234 280894 99854 298000
rect 100710 297805 100770 299510
rect 101446 297941 101506 299510
rect 101814 299510 101884 299570
rect 102912 299570 102972 300106
rect 103184 299842 103244 300106
rect 103184 299782 103346 299842
rect 102912 299510 102978 299570
rect 101814 298077 101874 299510
rect 102918 298213 102978 299510
rect 103286 298213 103346 299782
rect 104000 299570 104060 300106
rect 104408 299570 104468 300106
rect 105224 299842 105284 300106
rect 105224 299782 105370 299842
rect 104000 299510 104082 299570
rect 102915 298212 102981 298213
rect 102915 298148 102916 298212
rect 102980 298148 102981 298212
rect 102915 298147 102981 298148
rect 103283 298212 103349 298213
rect 103283 298148 103284 298212
rect 103348 298148 103349 298212
rect 103283 298147 103349 298148
rect 101811 298076 101877 298077
rect 101811 298012 101812 298076
rect 101876 298012 101877 298076
rect 101811 298011 101877 298012
rect 101443 297940 101509 297941
rect 101443 297876 101444 297940
rect 101508 297876 101509 297940
rect 101443 297875 101509 297876
rect 100707 297804 100773 297805
rect 100707 297740 100708 297804
rect 100772 297740 100773 297804
rect 100707 297739 100773 297740
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 132000 99854 136338
rect 102954 284614 103574 298000
rect 104022 297941 104082 299510
rect 104390 299510 104468 299570
rect 104390 298077 104450 299510
rect 104387 298076 104453 298077
rect 104387 298012 104388 298076
rect 104452 298012 104453 298076
rect 104387 298011 104453 298012
rect 105310 297941 105370 299782
rect 105632 299570 105692 300106
rect 106584 299570 106644 300106
rect 106856 299842 106916 300106
rect 106856 299782 107026 299842
rect 105632 299510 105738 299570
rect 106584 299510 106658 299570
rect 105678 298077 105738 299510
rect 106598 298077 106658 299510
rect 106966 298077 107026 299782
rect 107672 299570 107732 300106
rect 107808 299842 107868 300106
rect 107808 299782 107946 299842
rect 107672 299510 107762 299570
rect 105675 298076 105741 298077
rect 105675 298012 105676 298076
rect 105740 298012 105741 298076
rect 105675 298011 105741 298012
rect 106595 298076 106661 298077
rect 106595 298012 106596 298076
rect 106660 298012 106661 298076
rect 106595 298011 106661 298012
rect 106963 298076 107029 298077
rect 106963 298012 106964 298076
rect 107028 298012 107029 298076
rect 106963 298011 107029 298012
rect 107702 297941 107762 299510
rect 107886 298077 107946 299782
rect 109304 299570 109364 300106
rect 110528 299842 110588 300106
rect 110528 299782 110706 299842
rect 109304 299510 109418 299570
rect 109358 298077 109418 299510
rect 110646 298077 110706 299782
rect 111888 299570 111948 300106
rect 113112 299842 113172 300106
rect 113038 299782 113172 299842
rect 111888 299510 111994 299570
rect 107883 298076 107949 298077
rect 107883 298012 107884 298076
rect 107948 298012 107949 298076
rect 107883 298011 107949 298012
rect 109355 298076 109421 298077
rect 109355 298012 109356 298076
rect 109420 298012 109421 298076
rect 109355 298011 109421 298012
rect 110643 298076 110709 298077
rect 110643 298012 110644 298076
rect 110708 298012 110709 298076
rect 110643 298011 110709 298012
rect 104019 297940 104085 297941
rect 104019 297876 104020 297940
rect 104084 297876 104085 297940
rect 104019 297875 104085 297876
rect 105307 297940 105373 297941
rect 105307 297876 105308 297940
rect 105372 297876 105373 297940
rect 105307 297875 105373 297876
rect 107699 297940 107765 297941
rect 107699 297876 107700 297940
rect 107764 297876 107765 297940
rect 107699 297875 107765 297876
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 132000 103574 140058
rect 109794 291454 110414 298000
rect 111934 297941 111994 299510
rect 113038 298077 113098 299782
rect 114336 299570 114396 300106
rect 114326 299510 114396 299570
rect 115560 299570 115620 300106
rect 116784 299570 116844 300106
rect 115560 299510 115674 299570
rect 116784 299510 116962 299570
rect 114326 298077 114386 299510
rect 115614 298077 115674 299510
rect 116902 298077 116962 299510
rect 113035 298076 113101 298077
rect 113035 298012 113036 298076
rect 113100 298012 113101 298076
rect 113035 298011 113101 298012
rect 114323 298076 114389 298077
rect 114323 298012 114324 298076
rect 114388 298012 114389 298076
rect 114323 298011 114389 298012
rect 115611 298076 115677 298077
rect 115611 298012 115612 298076
rect 115676 298012 115677 298076
rect 115611 298011 115677 298012
rect 116899 298076 116965 298077
rect 116899 298012 116900 298076
rect 116964 298012 116965 298076
rect 116899 298011 116965 298012
rect 111931 297940 111997 297941
rect 111931 297876 111932 297940
rect 111996 297876 111997 297940
rect 111931 297875 111997 297876
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 132000 110414 146898
rect 113514 295174 114134 298000
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 132000 114134 150618
rect 117234 262894 117854 298000
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 132000 117854 154338
rect 120954 266614 121574 298000
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 132000 121574 158058
rect 127794 273454 128414 298000
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 132000 128414 164898
rect 131514 277174 132134 298000
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 132000 132134 132618
rect 135234 280894 135854 298000
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 34208 111454 34528 111486
rect 34208 111218 34250 111454
rect 34486 111218 34528 111454
rect 34208 111134 34528 111218
rect 34208 110898 34250 111134
rect 34486 110898 34528 111134
rect 34208 110866 34528 110898
rect 64928 111454 65248 111486
rect 64928 111218 64970 111454
rect 65206 111218 65248 111454
rect 64928 111134 65248 111218
rect 64928 110898 64970 111134
rect 65206 110898 65248 111134
rect 64928 110866 65248 110898
rect 95648 111454 95968 111486
rect 95648 111218 95690 111454
rect 95926 111218 95968 111454
rect 95648 111134 95968 111218
rect 95648 110898 95690 111134
rect 95926 110898 95968 111134
rect 95648 110866 95968 110898
rect 126368 111454 126688 111486
rect 126368 111218 126410 111454
rect 126646 111218 126688 111454
rect 126368 111134 126688 111218
rect 126368 110898 126410 111134
rect 126646 110898 126688 111134
rect 126368 110866 126688 110898
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 49568 93454 49888 93486
rect 49568 93218 49610 93454
rect 49846 93218 49888 93454
rect 49568 93134 49888 93218
rect 49568 92898 49610 93134
rect 49846 92898 49888 93134
rect 49568 92866 49888 92898
rect 80288 93454 80608 93486
rect 80288 93218 80330 93454
rect 80566 93218 80608 93454
rect 80288 93134 80608 93218
rect 80288 92898 80330 93134
rect 80566 92898 80608 93134
rect 80288 92866 80608 92898
rect 111008 93454 111328 93486
rect 111008 93218 111050 93454
rect 111286 93218 111328 93454
rect 111008 93134 111328 93218
rect 111008 92898 111050 93134
rect 111286 92898 111328 93134
rect 111008 92866 111328 92898
rect 34208 75454 34528 75486
rect 34208 75218 34250 75454
rect 34486 75218 34528 75454
rect 34208 75134 34528 75218
rect 34208 74898 34250 75134
rect 34486 74898 34528 75134
rect 34208 74866 34528 74898
rect 64928 75454 65248 75486
rect 64928 75218 64970 75454
rect 65206 75218 65248 75454
rect 64928 75134 65248 75218
rect 64928 74898 64970 75134
rect 65206 74898 65248 75134
rect 64928 74866 65248 74898
rect 95648 75454 95968 75486
rect 95648 75218 95690 75454
rect 95926 75218 95968 75454
rect 95648 75134 95968 75218
rect 95648 74898 95690 75134
rect 95926 74898 95968 75134
rect 95648 74866 95968 74898
rect 126368 75454 126688 75486
rect 126368 75218 126410 75454
rect 126646 75218 126688 75454
rect 126368 75134 126688 75218
rect 126368 74898 126410 75134
rect 126646 74898 126688 75134
rect 126368 74866 126688 74898
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 49568 57454 49888 57486
rect 49568 57218 49610 57454
rect 49846 57218 49888 57454
rect 49568 57134 49888 57218
rect 49568 56898 49610 57134
rect 49846 56898 49888 57134
rect 49568 56866 49888 56898
rect 80288 57454 80608 57486
rect 80288 57218 80330 57454
rect 80566 57218 80608 57454
rect 80288 57134 80608 57218
rect 80288 56898 80330 57134
rect 80566 56898 80608 57134
rect 80288 56866 80608 56898
rect 111008 57454 111328 57486
rect 111008 57218 111050 57454
rect 111286 57218 111328 57454
rect 111008 57134 111328 57218
rect 111008 56898 111050 57134
rect 111286 56898 111328 57134
rect 111008 56866 111328 56898
rect 34208 39454 34528 39486
rect 34208 39218 34250 39454
rect 34486 39218 34528 39454
rect 34208 39134 34528 39218
rect 34208 38898 34250 39134
rect 34486 38898 34528 39134
rect 34208 38866 34528 38898
rect 64928 39454 65248 39486
rect 64928 39218 64970 39454
rect 65206 39218 65248 39454
rect 64928 39134 65248 39218
rect 64928 38898 64970 39134
rect 65206 38898 65248 39134
rect 64928 38866 65248 38898
rect 95648 39454 95968 39486
rect 95648 39218 95690 39454
rect 95926 39218 95968 39454
rect 95648 39134 95968 39218
rect 95648 38898 95690 39134
rect 95926 38898 95968 39134
rect 95648 38866 95968 38898
rect 126368 39454 126688 39486
rect 126368 39218 126410 39454
rect 126646 39218 126688 39454
rect 126368 39134 126688 39218
rect 126368 38898 126410 39134
rect 126646 38898 126688 39134
rect 126368 38866 126688 38898
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 28000
rect 37794 3454 38414 28000
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 7174 42134 28000
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 10894 45854 28000
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 14614 49574 28000
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 28000
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 28000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 28000
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 28000
rect 73794 3454 74414 28000
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 7174 78134 28000
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 10894 81854 28000
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 14614 85574 28000
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 21454 92414 28000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 28000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 -5146 99854 28000
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 28000
rect 109794 3454 110414 28000
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 7174 114134 28000
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 10894 117854 28000
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 14614 121574 28000
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 21454 128414 28000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 28000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 284614 139574 298000
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 291454 146414 298000
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 252000 189854 262338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 252000 193574 266058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 252000 200414 272898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 252000 204134 276618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 381500 211574 392058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 381500 218414 398898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 381500 222134 402618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 381500 225854 406338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 381500 229574 410058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381500 236414 416898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 381500 240134 384618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 381500 243854 388338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 381500 247574 392058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 381500 254414 398898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 381500 258134 402618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 381500 261854 406338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 381500 265574 410058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381500 272414 416898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 381500 276134 384618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 381500 279854 388338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 381500 283574 392058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 381500 290414 398898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 381500 294134 402618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 381500 297854 406338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 381500 301574 410058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381500 308414 416898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 210952 363454 211300 363486
rect 210952 363218 211008 363454
rect 211244 363218 211300 363454
rect 210952 363134 211300 363218
rect 210952 362898 211008 363134
rect 211244 362898 211300 363134
rect 210952 362866 211300 362898
rect 304656 363454 305004 363486
rect 304656 363218 304712 363454
rect 304948 363218 305004 363454
rect 304656 363134 305004 363218
rect 304656 362898 304712 363134
rect 304948 362898 305004 363134
rect 304656 362866 305004 362898
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 210272 345454 210620 345486
rect 210272 345218 210328 345454
rect 210564 345218 210620 345454
rect 210272 345134 210620 345218
rect 210272 344898 210328 345134
rect 210564 344898 210620 345134
rect 210272 344866 210620 344898
rect 305336 345454 305684 345486
rect 305336 345218 305392 345454
rect 305628 345218 305684 345454
rect 305336 345134 305684 345218
rect 305336 344898 305392 345134
rect 305628 344898 305684 345134
rect 305336 344866 305684 344898
rect 210952 327454 211300 327486
rect 210952 327218 211008 327454
rect 211244 327218 211300 327454
rect 210952 327134 211300 327218
rect 210952 326898 211008 327134
rect 211244 326898 211300 327134
rect 210952 326866 211300 326898
rect 304656 327454 305004 327486
rect 304656 327218 304712 327454
rect 304948 327218 305004 327454
rect 304656 327134 305004 327218
rect 304656 326898 304712 327134
rect 304948 326898 305004 327134
rect 304656 326866 305004 326898
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 210272 309454 210620 309486
rect 210272 309218 210328 309454
rect 210564 309218 210620 309454
rect 210272 309134 210620 309218
rect 210272 308898 210328 309134
rect 210564 308898 210620 309134
rect 210272 308866 210620 308898
rect 305336 309454 305684 309486
rect 305336 309218 305392 309454
rect 305628 309218 305684 309454
rect 305336 309134 305684 309218
rect 305336 308898 305392 309134
rect 305628 308898 305684 309134
rect 305336 308866 305684 308898
rect 215856 299570 215916 300106
rect 225512 299570 225572 300106
rect 215856 299510 215954 299570
rect 215894 298077 215954 299510
rect 225462 299510 225572 299570
rect 226736 299570 226796 300106
rect 227824 299570 227884 300106
rect 229184 299570 229244 300106
rect 230136 299570 230196 300106
rect 231360 299570 231420 300106
rect 226736 299510 226810 299570
rect 227824 299510 227914 299570
rect 225462 298213 225522 299510
rect 225459 298212 225525 298213
rect 225459 298148 225460 298212
rect 225524 298148 225525 298212
rect 225459 298147 225525 298148
rect 226750 298077 226810 299510
rect 227854 298077 227914 299510
rect 229142 299510 229244 299570
rect 230062 299510 230196 299570
rect 231350 299510 231420 299570
rect 232584 299570 232644 300106
rect 233672 299570 233732 300106
rect 235032 299570 235092 300106
rect 232584 299510 232698 299570
rect 229142 298213 229202 299510
rect 229139 298212 229205 298213
rect 229139 298148 229140 298212
rect 229204 298148 229205 298212
rect 229139 298147 229205 298148
rect 215891 298076 215957 298077
rect 215891 298012 215892 298076
rect 215956 298012 215957 298076
rect 215891 298011 215957 298012
rect 226747 298076 226813 298077
rect 226747 298012 226748 298076
rect 226812 298012 226813 298076
rect 226747 298011 226813 298012
rect 227851 298076 227917 298077
rect 227851 298012 227852 298076
rect 227916 298012 227917 298076
rect 227851 298011 227917 298012
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 252000 207854 280338
rect 210954 284614 211574 298000
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 252000 211574 284058
rect 217794 291454 218414 298000
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 252000 218414 254898
rect 221514 295174 222134 298000
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 252000 222134 258618
rect 225234 262894 225854 298000
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 252000 225854 262338
rect 228954 266614 229574 298000
rect 230062 297261 230122 299510
rect 231350 298077 231410 299510
rect 232638 298077 232698 299510
rect 233558 299510 233732 299570
rect 235030 299510 235092 299570
rect 236120 299570 236180 300106
rect 237208 299570 237268 300106
rect 237888 299570 237948 300106
rect 236120 299510 236562 299570
rect 237208 299510 237298 299570
rect 233558 298077 233618 299510
rect 235030 298077 235090 299510
rect 231347 298076 231413 298077
rect 231347 298012 231348 298076
rect 231412 298012 231413 298076
rect 231347 298011 231413 298012
rect 232635 298076 232701 298077
rect 232635 298012 232636 298076
rect 232700 298012 232701 298076
rect 232635 298011 232701 298012
rect 233555 298076 233621 298077
rect 233555 298012 233556 298076
rect 233620 298012 233621 298076
rect 233555 298011 233621 298012
rect 235027 298076 235093 298077
rect 235027 298012 235028 298076
rect 235092 298012 235093 298076
rect 235027 298011 235093 298012
rect 230059 297260 230125 297261
rect 230059 297196 230060 297260
rect 230124 297196 230125 297260
rect 230059 297195 230125 297196
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 252000 229574 266058
rect 235794 273454 236414 298000
rect 236502 297805 236562 299510
rect 237238 298077 237298 299510
rect 237790 299510 237948 299570
rect 238296 299570 238356 300106
rect 239248 299570 239308 300106
rect 239656 299845 239716 300106
rect 239653 299844 239719 299845
rect 239653 299780 239654 299844
rect 239718 299780 239719 299844
rect 239653 299779 239719 299780
rect 240336 299570 240396 300106
rect 240744 299570 240804 300106
rect 238296 299510 238402 299570
rect 239248 299510 239322 299570
rect 240336 299510 240426 299570
rect 237235 298076 237301 298077
rect 237235 298012 237236 298076
rect 237300 298012 237301 298076
rect 237235 298011 237301 298012
rect 237790 297941 237850 299510
rect 237787 297940 237853 297941
rect 237787 297876 237788 297940
rect 237852 297876 237853 297940
rect 237787 297875 237853 297876
rect 236499 297804 236565 297805
rect 236499 297740 236500 297804
rect 236564 297740 236565 297804
rect 236499 297739 236565 297740
rect 238342 296853 238402 299510
rect 239262 298077 239322 299510
rect 240366 298077 240426 299510
rect 240734 299510 240804 299570
rect 241832 299570 241892 300106
rect 241968 299570 242028 300106
rect 243056 299709 243116 300106
rect 243053 299708 243119 299709
rect 243053 299644 243054 299708
rect 243118 299644 243119 299708
rect 243053 299643 243119 299644
rect 243192 299570 243252 300106
rect 244144 299570 244204 300106
rect 244416 299570 244476 300106
rect 241832 299510 241898 299570
rect 241968 299510 242082 299570
rect 240734 298077 240794 299510
rect 239259 298076 239325 298077
rect 239259 298012 239260 298076
rect 239324 298012 239325 298076
rect 239259 298011 239325 298012
rect 240363 298076 240429 298077
rect 240363 298012 240364 298076
rect 240428 298012 240429 298076
rect 240363 298011 240429 298012
rect 240731 298076 240797 298077
rect 240731 298012 240732 298076
rect 240796 298012 240797 298076
rect 240731 298011 240797 298012
rect 238339 296852 238405 296853
rect 238339 296788 238340 296852
rect 238404 296788 238405 296852
rect 238339 296787 238405 296788
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 252000 236414 272898
rect 239514 277174 240134 298000
rect 241838 297805 241898 299510
rect 242022 297941 242082 299510
rect 242942 299510 243252 299570
rect 244046 299510 244204 299570
rect 244414 299510 244476 299570
rect 245504 299570 245564 300106
rect 245640 299570 245700 300106
rect 246592 299570 246652 300106
rect 246864 299570 246924 300106
rect 247680 299570 247740 300106
rect 245504 299510 245578 299570
rect 245640 299510 245762 299570
rect 246592 299510 246682 299570
rect 242942 298077 243002 299510
rect 244046 298077 244106 299510
rect 244414 298077 244474 299510
rect 245518 298077 245578 299510
rect 242939 298076 243005 298077
rect 242939 298012 242940 298076
rect 243004 298012 243005 298076
rect 242939 298011 243005 298012
rect 244043 298076 244109 298077
rect 244043 298012 244044 298076
rect 244108 298012 244109 298076
rect 244043 298011 244109 298012
rect 244411 298076 244477 298077
rect 244411 298012 244412 298076
rect 244476 298012 244477 298076
rect 244411 298011 244477 298012
rect 245515 298076 245581 298077
rect 245515 298012 245516 298076
rect 245580 298012 245581 298076
rect 245515 298011 245581 298012
rect 242019 297940 242085 297941
rect 242019 297876 242020 297940
rect 242084 297876 242085 297940
rect 242019 297875 242085 297876
rect 241835 297804 241901 297805
rect 241835 297740 241836 297804
rect 241900 297740 241901 297804
rect 241835 297739 241901 297740
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 252000 240134 276618
rect 243234 280894 243854 298000
rect 245702 297805 245762 299510
rect 246622 297941 246682 299510
rect 246806 299510 246924 299570
rect 247542 299510 247740 299570
rect 247816 299570 247876 300106
rect 248904 299842 248964 300106
rect 249312 299842 249372 300106
rect 248904 299782 249074 299842
rect 249312 299782 249442 299842
rect 247816 299510 247970 299570
rect 246806 298077 246866 299510
rect 247542 298890 247602 299510
rect 247542 298830 247786 298890
rect 246803 298076 246869 298077
rect 246803 298012 246804 298076
rect 246868 298012 246869 298076
rect 246803 298011 246869 298012
rect 246619 297940 246685 297941
rect 246619 297876 246620 297940
rect 246684 297876 246685 297940
rect 246619 297875 246685 297876
rect 245699 297804 245765 297805
rect 245699 297740 245700 297804
rect 245764 297740 245765 297804
rect 245699 297739 245765 297740
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 252000 243854 280338
rect 246954 284614 247574 298000
rect 247726 297941 247786 298830
rect 247910 298077 247970 299510
rect 247907 298076 247973 298077
rect 247907 298012 247908 298076
rect 247972 298012 247973 298076
rect 247907 298011 247973 298012
rect 249014 297941 249074 299782
rect 249382 298077 249442 299782
rect 250264 299570 250324 300106
rect 250672 299570 250732 300106
rect 250264 299510 250362 299570
rect 249379 298076 249445 298077
rect 249379 298012 249380 298076
rect 249444 298012 249445 298076
rect 249379 298011 249445 298012
rect 250302 297941 250362 299510
rect 250670 299510 250732 299570
rect 251352 299570 251412 300106
rect 251896 299570 251956 300106
rect 252440 299842 252500 300106
rect 252440 299782 252570 299842
rect 251352 299510 251466 299570
rect 251896 299510 252018 299570
rect 250670 298077 250730 299510
rect 250667 298076 250733 298077
rect 250667 298012 250668 298076
rect 250732 298012 250733 298076
rect 250667 298011 250733 298012
rect 251406 297941 251466 299510
rect 247723 297940 247789 297941
rect 247723 297876 247724 297940
rect 247788 297876 247789 297940
rect 247723 297875 247789 297876
rect 249011 297940 249077 297941
rect 249011 297876 249012 297940
rect 249076 297876 249077 297940
rect 249011 297875 249077 297876
rect 250299 297940 250365 297941
rect 250299 297876 250300 297940
rect 250364 297876 250365 297940
rect 250299 297875 250365 297876
rect 251403 297940 251469 297941
rect 251403 297876 251404 297940
rect 251468 297876 251469 297940
rect 251403 297875 251469 297876
rect 251958 297805 252018 299510
rect 252510 298077 252570 299782
rect 253120 299570 253180 300106
rect 253528 299842 253588 300106
rect 253528 299782 253674 299842
rect 253062 299510 253180 299570
rect 252507 298076 252573 298077
rect 252507 298012 252508 298076
rect 252572 298012 252573 298076
rect 252507 298011 252573 298012
rect 253062 297941 253122 299510
rect 253614 298077 253674 299782
rect 254344 299570 254404 300106
rect 254888 299570 254948 300106
rect 255568 299842 255628 300106
rect 255568 299782 255698 299842
rect 254344 299510 254594 299570
rect 254888 299510 254962 299570
rect 253611 298076 253677 298077
rect 253611 298012 253612 298076
rect 253676 298012 253677 298076
rect 253611 298011 253677 298012
rect 253059 297940 253125 297941
rect 253059 297876 253060 297940
rect 253124 297876 253125 297940
rect 253059 297875 253125 297876
rect 251955 297804 252021 297805
rect 251955 297740 251956 297804
rect 252020 297740 252021 297804
rect 251955 297739 252021 297740
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 252000 247574 284058
rect 253794 291454 254414 298000
rect 254534 297941 254594 299510
rect 254902 298077 254962 299510
rect 254899 298076 254965 298077
rect 254899 298012 254900 298076
rect 254964 298012 254965 298076
rect 254899 298011 254965 298012
rect 255638 297941 255698 299782
rect 255976 299570 256036 300106
rect 256656 299842 256716 300106
rect 256656 299782 256802 299842
rect 255976 299510 256066 299570
rect 256006 298077 256066 299510
rect 256003 298076 256069 298077
rect 256003 298012 256004 298076
rect 256068 298012 256069 298076
rect 256003 298011 256069 298012
rect 256742 297941 256802 299782
rect 257064 299570 257124 300106
rect 257880 299570 257940 300106
rect 257064 299510 257170 299570
rect 257110 298077 257170 299510
rect 257846 299510 257940 299570
rect 258288 299570 258348 300106
rect 259104 299570 259164 300106
rect 259376 299570 259436 300106
rect 258288 299510 258458 299570
rect 259104 299510 259194 299570
rect 257846 298213 257906 299510
rect 257843 298212 257909 298213
rect 257843 298148 257844 298212
rect 257908 298148 257909 298212
rect 257843 298147 257909 298148
rect 257107 298076 257173 298077
rect 257107 298012 257108 298076
rect 257172 298012 257173 298076
rect 257107 298011 257173 298012
rect 254531 297940 254597 297941
rect 254531 297876 254532 297940
rect 254596 297876 254597 297940
rect 254531 297875 254597 297876
rect 255635 297940 255701 297941
rect 255635 297876 255636 297940
rect 255700 297876 255701 297940
rect 255635 297875 255701 297876
rect 256739 297940 256805 297941
rect 256739 297876 256740 297940
rect 256804 297876 256805 297940
rect 256739 297875 256805 297876
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 252000 254414 254898
rect 257514 295174 258134 298000
rect 258398 297805 258458 299510
rect 259134 297941 259194 299510
rect 259318 299510 259436 299570
rect 260600 299570 260660 300106
rect 260736 299570 260796 300106
rect 261416 299570 261476 300106
rect 261824 299570 261884 300106
rect 262912 299570 262972 300106
rect 263184 299570 263244 300106
rect 260600 299510 260666 299570
rect 260736 299510 260850 299570
rect 261416 299510 261586 299570
rect 261824 299510 261954 299570
rect 262912 299510 263058 299570
rect 259318 298077 259378 299510
rect 259315 298076 259381 298077
rect 259315 298012 259316 298076
rect 259380 298012 259381 298076
rect 259315 298011 259381 298012
rect 260606 297941 260666 299510
rect 260790 298077 260850 299510
rect 261526 298213 261586 299510
rect 261894 298213 261954 299510
rect 261523 298212 261589 298213
rect 261523 298148 261524 298212
rect 261588 298148 261589 298212
rect 261523 298147 261589 298148
rect 261891 298212 261957 298213
rect 261891 298148 261892 298212
rect 261956 298148 261957 298212
rect 261891 298147 261957 298148
rect 260787 298076 260853 298077
rect 260787 298012 260788 298076
rect 260852 298012 260853 298076
rect 260787 298011 260853 298012
rect 259131 297940 259197 297941
rect 259131 297876 259132 297940
rect 259196 297876 259197 297940
rect 259131 297875 259197 297876
rect 260603 297940 260669 297941
rect 260603 297876 260604 297940
rect 260668 297876 260669 297940
rect 260603 297875 260669 297876
rect 258395 297804 258461 297805
rect 258395 297740 258396 297804
rect 258460 297740 258461 297804
rect 258395 297739 258461 297740
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 252000 258134 258618
rect 261234 262894 261854 298000
rect 262998 297941 263058 299510
rect 263182 299510 263244 299570
rect 264000 299570 264060 300106
rect 264408 299570 264468 300106
rect 265224 299570 265284 300106
rect 264000 299510 264162 299570
rect 264408 299510 264530 299570
rect 263182 298077 263242 299510
rect 263179 298076 263245 298077
rect 263179 298012 263180 298076
rect 263244 298012 263245 298076
rect 263179 298011 263245 298012
rect 262995 297940 263061 297941
rect 262995 297876 262996 297940
rect 263060 297876 263061 297940
rect 262995 297875 263061 297876
rect 264102 296989 264162 299510
rect 264099 296988 264165 296989
rect 264099 296924 264100 296988
rect 264164 296924 264165 296988
rect 264099 296923 264165 296924
rect 264470 296853 264530 299510
rect 265206 299510 265284 299570
rect 265632 299570 265692 300106
rect 266584 299570 266644 300106
rect 266856 299570 266916 300106
rect 267672 299570 267732 300106
rect 265632 299510 265818 299570
rect 266584 299510 266738 299570
rect 266856 299510 266922 299570
rect 265206 298213 265266 299510
rect 265203 298212 265269 298213
rect 265203 298148 265204 298212
rect 265268 298148 265269 298212
rect 265203 298147 265269 298148
rect 264467 296852 264533 296853
rect 264467 296788 264468 296852
rect 264532 296788 264533 296852
rect 264467 296787 264533 296788
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 252000 261854 262338
rect 264954 266614 265574 298000
rect 265758 296853 265818 299510
rect 266678 297125 266738 299510
rect 266675 297124 266741 297125
rect 266675 297060 266676 297124
rect 266740 297060 266741 297124
rect 266675 297059 266741 297060
rect 266862 296989 266922 299510
rect 267598 299510 267732 299570
rect 267808 299570 267868 300106
rect 269304 299570 269364 300106
rect 267808 299510 268026 299570
rect 266859 296988 266925 296989
rect 266859 296924 266860 296988
rect 266924 296924 266925 296988
rect 266859 296923 266925 296924
rect 267598 296853 267658 299510
rect 267966 297533 268026 299510
rect 269254 299510 269364 299570
rect 270528 299570 270588 300106
rect 271888 299570 271948 300106
rect 270528 299510 270602 299570
rect 267963 297532 268029 297533
rect 267963 297468 267964 297532
rect 268028 297468 268029 297532
rect 267963 297467 268029 297468
rect 269254 296853 269314 299510
rect 270542 296853 270602 299510
rect 271830 299510 271948 299570
rect 273112 299570 273172 300106
rect 274336 299842 274396 300106
rect 274336 299782 274466 299842
rect 273112 299510 273178 299570
rect 271830 298213 271890 299510
rect 271827 298212 271893 298213
rect 271827 298148 271828 298212
rect 271892 298148 271893 298212
rect 271827 298147 271893 298148
rect 265755 296852 265821 296853
rect 265755 296788 265756 296852
rect 265820 296788 265821 296852
rect 265755 296787 265821 296788
rect 267595 296852 267661 296853
rect 267595 296788 267596 296852
rect 267660 296788 267661 296852
rect 267595 296787 267661 296788
rect 269251 296852 269317 296853
rect 269251 296788 269252 296852
rect 269316 296788 269317 296852
rect 269251 296787 269317 296788
rect 270539 296852 270605 296853
rect 270539 296788 270540 296852
rect 270604 296788 270605 296852
rect 270539 296787 270605 296788
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 252000 265574 266058
rect 271794 273454 272414 298000
rect 273118 296853 273178 299510
rect 274406 298077 274466 299782
rect 275560 299570 275620 300106
rect 275510 299510 275620 299570
rect 276784 299570 276844 300106
rect 276784 299510 276858 299570
rect 275510 298213 275570 299510
rect 275507 298212 275573 298213
rect 275507 298148 275508 298212
rect 275572 298148 275573 298212
rect 275507 298147 275573 298148
rect 276798 298077 276858 299510
rect 274403 298076 274469 298077
rect 274403 298012 274404 298076
rect 274468 298012 274469 298076
rect 274403 298011 274469 298012
rect 276795 298076 276861 298077
rect 276795 298012 276796 298076
rect 276860 298012 276861 298076
rect 276795 298011 276861 298012
rect 273115 296852 273181 296853
rect 273115 296788 273116 296852
rect 273180 296788 273181 296852
rect 273115 296787 273181 296788
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 252000 272414 272898
rect 275514 277174 276134 298000
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 252000 276134 276618
rect 279234 280894 279854 298000
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 252000 279854 280338
rect 282954 284614 283574 298000
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 252000 283574 284058
rect 289794 291454 290414 298000
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 252000 290414 254898
rect 293514 295174 294134 298000
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 252000 294134 258618
rect 297234 262894 297854 298000
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 252000 297854 262338
rect 300954 266614 301574 298000
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 252000 301574 266058
rect 307794 273454 308414 298000
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 252000 308414 272898
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 252000 312134 276618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 252000 315854 280338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 252000 319574 284058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 252000 326414 254898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 252000 330134 258618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 252000 333854 262338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 252000 337574 266058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 252000 344414 272898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 252000 348134 276618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 252000 351854 280338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 252000 355574 284058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 252000 362414 254898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 252000 366134 258618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 252000 369854 262338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 252000 373574 266058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 252000 380414 272898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 252000 384134 276618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 252000 387854 280338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 252000 391574 284058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 252000 398414 254898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 252000 402134 258618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 252000 405854 262338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 252000 409574 266058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 209568 237454 209888 237486
rect 209568 237218 209610 237454
rect 209846 237218 209888 237454
rect 209568 237134 209888 237218
rect 209568 236898 209610 237134
rect 209846 236898 209888 237134
rect 209568 236866 209888 236898
rect 240288 237454 240608 237486
rect 240288 237218 240330 237454
rect 240566 237218 240608 237454
rect 240288 237134 240608 237218
rect 240288 236898 240330 237134
rect 240566 236898 240608 237134
rect 240288 236866 240608 236898
rect 271008 237454 271328 237486
rect 271008 237218 271050 237454
rect 271286 237218 271328 237454
rect 271008 237134 271328 237218
rect 271008 236898 271050 237134
rect 271286 236898 271328 237134
rect 271008 236866 271328 236898
rect 301728 237454 302048 237486
rect 301728 237218 301770 237454
rect 302006 237218 302048 237454
rect 301728 237134 302048 237218
rect 301728 236898 301770 237134
rect 302006 236898 302048 237134
rect 301728 236866 302048 236898
rect 332448 237454 332768 237486
rect 332448 237218 332490 237454
rect 332726 237218 332768 237454
rect 332448 237134 332768 237218
rect 332448 236898 332490 237134
rect 332726 236898 332768 237134
rect 332448 236866 332768 236898
rect 363168 237454 363488 237486
rect 363168 237218 363210 237454
rect 363446 237218 363488 237454
rect 363168 237134 363488 237218
rect 363168 236898 363210 237134
rect 363446 236898 363488 237134
rect 363168 236866 363488 236898
rect 393888 237454 394208 237486
rect 393888 237218 393930 237454
rect 394166 237218 394208 237454
rect 393888 237134 394208 237218
rect 393888 236898 393930 237134
rect 394166 236898 394208 237134
rect 393888 236866 394208 236898
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 194208 219454 194528 219486
rect 194208 219218 194250 219454
rect 194486 219218 194528 219454
rect 194208 219134 194528 219218
rect 194208 218898 194250 219134
rect 194486 218898 194528 219134
rect 194208 218866 194528 218898
rect 224928 219454 225248 219486
rect 224928 219218 224970 219454
rect 225206 219218 225248 219454
rect 224928 219134 225248 219218
rect 224928 218898 224970 219134
rect 225206 218898 225248 219134
rect 224928 218866 225248 218898
rect 255648 219454 255968 219486
rect 255648 219218 255690 219454
rect 255926 219218 255968 219454
rect 255648 219134 255968 219218
rect 255648 218898 255690 219134
rect 255926 218898 255968 219134
rect 255648 218866 255968 218898
rect 286368 219454 286688 219486
rect 286368 219218 286410 219454
rect 286646 219218 286688 219454
rect 286368 219134 286688 219218
rect 286368 218898 286410 219134
rect 286646 218898 286688 219134
rect 286368 218866 286688 218898
rect 317088 219454 317408 219486
rect 317088 219218 317130 219454
rect 317366 219218 317408 219454
rect 317088 219134 317408 219218
rect 317088 218898 317130 219134
rect 317366 218898 317408 219134
rect 317088 218866 317408 218898
rect 347808 219454 348128 219486
rect 347808 219218 347850 219454
rect 348086 219218 348128 219454
rect 347808 219134 348128 219218
rect 347808 218898 347850 219134
rect 348086 218898 348128 219134
rect 347808 218866 348128 218898
rect 378528 219454 378848 219486
rect 378528 219218 378570 219454
rect 378806 219218 378848 219454
rect 378528 219134 378848 219218
rect 378528 218898 378570 219134
rect 378806 218898 378848 219134
rect 378528 218866 378848 218898
rect 209568 201454 209888 201486
rect 209568 201218 209610 201454
rect 209846 201218 209888 201454
rect 209568 201134 209888 201218
rect 209568 200898 209610 201134
rect 209846 200898 209888 201134
rect 209568 200866 209888 200898
rect 240288 201454 240608 201486
rect 240288 201218 240330 201454
rect 240566 201218 240608 201454
rect 240288 201134 240608 201218
rect 240288 200898 240330 201134
rect 240566 200898 240608 201134
rect 240288 200866 240608 200898
rect 271008 201454 271328 201486
rect 271008 201218 271050 201454
rect 271286 201218 271328 201454
rect 271008 201134 271328 201218
rect 271008 200898 271050 201134
rect 271286 200898 271328 201134
rect 271008 200866 271328 200898
rect 301728 201454 302048 201486
rect 301728 201218 301770 201454
rect 302006 201218 302048 201454
rect 301728 201134 302048 201218
rect 301728 200898 301770 201134
rect 302006 200898 302048 201134
rect 301728 200866 302048 200898
rect 332448 201454 332768 201486
rect 332448 201218 332490 201454
rect 332726 201218 332768 201454
rect 332448 201134 332768 201218
rect 332448 200898 332490 201134
rect 332726 200898 332768 201134
rect 332448 200866 332768 200898
rect 363168 201454 363488 201486
rect 363168 201218 363210 201454
rect 363446 201218 363488 201454
rect 363168 201134 363488 201218
rect 363168 200898 363210 201134
rect 363446 200898 363488 201134
rect 363168 200866 363488 200898
rect 393888 201454 394208 201486
rect 393888 201218 393930 201454
rect 394166 201218 394208 201454
rect 393888 201134 394208 201218
rect 393888 200898 393930 201134
rect 394166 200898 394208 201134
rect 393888 200866 394208 200898
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 194208 183454 194528 183486
rect 194208 183218 194250 183454
rect 194486 183218 194528 183454
rect 194208 183134 194528 183218
rect 194208 182898 194250 183134
rect 194486 182898 194528 183134
rect 194208 182866 194528 182898
rect 224928 183454 225248 183486
rect 224928 183218 224970 183454
rect 225206 183218 225248 183454
rect 224928 183134 225248 183218
rect 224928 182898 224970 183134
rect 225206 182898 225248 183134
rect 224928 182866 225248 182898
rect 255648 183454 255968 183486
rect 255648 183218 255690 183454
rect 255926 183218 255968 183454
rect 255648 183134 255968 183218
rect 255648 182898 255690 183134
rect 255926 182898 255968 183134
rect 255648 182866 255968 182898
rect 286368 183454 286688 183486
rect 286368 183218 286410 183454
rect 286646 183218 286688 183454
rect 286368 183134 286688 183218
rect 286368 182898 286410 183134
rect 286646 182898 286688 183134
rect 286368 182866 286688 182898
rect 317088 183454 317408 183486
rect 317088 183218 317130 183454
rect 317366 183218 317408 183454
rect 317088 183134 317408 183218
rect 317088 182898 317130 183134
rect 317366 182898 317408 183134
rect 317088 182866 317408 182898
rect 347808 183454 348128 183486
rect 347808 183218 347850 183454
rect 348086 183218 348128 183454
rect 347808 183134 348128 183218
rect 347808 182898 347850 183134
rect 348086 182898 348128 183134
rect 347808 182866 348128 182898
rect 378528 183454 378848 183486
rect 378528 183218 378570 183454
rect 378806 183218 378848 183454
rect 378528 183134 378848 183218
rect 378528 182898 378570 183134
rect 378806 182898 378848 183134
rect 378528 182866 378848 182898
rect 209568 165454 209888 165486
rect 209568 165218 209610 165454
rect 209846 165218 209888 165454
rect 209568 165134 209888 165218
rect 209568 164898 209610 165134
rect 209846 164898 209888 165134
rect 209568 164866 209888 164898
rect 240288 165454 240608 165486
rect 240288 165218 240330 165454
rect 240566 165218 240608 165454
rect 240288 165134 240608 165218
rect 240288 164898 240330 165134
rect 240566 164898 240608 165134
rect 240288 164866 240608 164898
rect 271008 165454 271328 165486
rect 271008 165218 271050 165454
rect 271286 165218 271328 165454
rect 271008 165134 271328 165218
rect 271008 164898 271050 165134
rect 271286 164898 271328 165134
rect 271008 164866 271328 164898
rect 301728 165454 302048 165486
rect 301728 165218 301770 165454
rect 302006 165218 302048 165454
rect 301728 165134 302048 165218
rect 301728 164898 301770 165134
rect 302006 164898 302048 165134
rect 301728 164866 302048 164898
rect 332448 165454 332768 165486
rect 332448 165218 332490 165454
rect 332726 165218 332768 165454
rect 332448 165134 332768 165218
rect 332448 164898 332490 165134
rect 332726 164898 332768 165134
rect 332448 164866 332768 164898
rect 363168 165454 363488 165486
rect 363168 165218 363210 165454
rect 363446 165218 363488 165454
rect 363168 165134 363488 165218
rect 363168 164898 363210 165134
rect 363446 164898 363488 165134
rect 363168 164866 363488 164898
rect 393888 165454 394208 165486
rect 393888 165218 393930 165454
rect 394166 165218 394208 165454
rect 393888 165134 394208 165218
rect 393888 164898 393930 165134
rect 394166 164898 394208 165134
rect 393888 164866 394208 164898
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 194208 147454 194528 147486
rect 194208 147218 194250 147454
rect 194486 147218 194528 147454
rect 194208 147134 194528 147218
rect 194208 146898 194250 147134
rect 194486 146898 194528 147134
rect 194208 146866 194528 146898
rect 224928 147454 225248 147486
rect 224928 147218 224970 147454
rect 225206 147218 225248 147454
rect 224928 147134 225248 147218
rect 224928 146898 224970 147134
rect 225206 146898 225248 147134
rect 224928 146866 225248 146898
rect 255648 147454 255968 147486
rect 255648 147218 255690 147454
rect 255926 147218 255968 147454
rect 255648 147134 255968 147218
rect 255648 146898 255690 147134
rect 255926 146898 255968 147134
rect 255648 146866 255968 146898
rect 286368 147454 286688 147486
rect 286368 147218 286410 147454
rect 286646 147218 286688 147454
rect 286368 147134 286688 147218
rect 286368 146898 286410 147134
rect 286646 146898 286688 147134
rect 286368 146866 286688 146898
rect 317088 147454 317408 147486
rect 317088 147218 317130 147454
rect 317366 147218 317408 147454
rect 317088 147134 317408 147218
rect 317088 146898 317130 147134
rect 317366 146898 317408 147134
rect 317088 146866 317408 146898
rect 347808 147454 348128 147486
rect 347808 147218 347850 147454
rect 348086 147218 348128 147454
rect 347808 147134 348128 147218
rect 347808 146898 347850 147134
rect 348086 146898 348128 147134
rect 347808 146866 348128 146898
rect 378528 147454 378848 147486
rect 378528 147218 378570 147454
rect 378806 147218 378848 147454
rect 378528 147134 378848 147218
rect 378528 146898 378570 147134
rect 378806 146898 378848 147134
rect 378528 146866 378848 146898
rect 209568 129454 209888 129486
rect 209568 129218 209610 129454
rect 209846 129218 209888 129454
rect 209568 129134 209888 129218
rect 209568 128898 209610 129134
rect 209846 128898 209888 129134
rect 209568 128866 209888 128898
rect 240288 129454 240608 129486
rect 240288 129218 240330 129454
rect 240566 129218 240608 129454
rect 240288 129134 240608 129218
rect 240288 128898 240330 129134
rect 240566 128898 240608 129134
rect 240288 128866 240608 128898
rect 271008 129454 271328 129486
rect 271008 129218 271050 129454
rect 271286 129218 271328 129454
rect 271008 129134 271328 129218
rect 271008 128898 271050 129134
rect 271286 128898 271328 129134
rect 271008 128866 271328 128898
rect 301728 129454 302048 129486
rect 301728 129218 301770 129454
rect 302006 129218 302048 129454
rect 301728 129134 302048 129218
rect 301728 128898 301770 129134
rect 302006 128898 302048 129134
rect 301728 128866 302048 128898
rect 332448 129454 332768 129486
rect 332448 129218 332490 129454
rect 332726 129218 332768 129454
rect 332448 129134 332768 129218
rect 332448 128898 332490 129134
rect 332726 128898 332768 129134
rect 332448 128866 332768 128898
rect 363168 129454 363488 129486
rect 363168 129218 363210 129454
rect 363446 129218 363488 129454
rect 363168 129134 363488 129218
rect 363168 128898 363210 129134
rect 363446 128898 363488 129134
rect 363168 128866 363488 128898
rect 393888 129454 394208 129486
rect 393888 129218 393930 129454
rect 394166 129218 394208 129454
rect 393888 129134 394208 129218
rect 393888 128898 393930 129134
rect 394166 128898 394208 129134
rect 393888 128866 394208 128898
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 194208 111454 194528 111486
rect 194208 111218 194250 111454
rect 194486 111218 194528 111454
rect 194208 111134 194528 111218
rect 194208 110898 194250 111134
rect 194486 110898 194528 111134
rect 194208 110866 194528 110898
rect 224928 111454 225248 111486
rect 224928 111218 224970 111454
rect 225206 111218 225248 111454
rect 224928 111134 225248 111218
rect 224928 110898 224970 111134
rect 225206 110898 225248 111134
rect 224928 110866 225248 110898
rect 255648 111454 255968 111486
rect 255648 111218 255690 111454
rect 255926 111218 255968 111454
rect 255648 111134 255968 111218
rect 255648 110898 255690 111134
rect 255926 110898 255968 111134
rect 255648 110866 255968 110898
rect 286368 111454 286688 111486
rect 286368 111218 286410 111454
rect 286646 111218 286688 111454
rect 286368 111134 286688 111218
rect 286368 110898 286410 111134
rect 286646 110898 286688 111134
rect 286368 110866 286688 110898
rect 317088 111454 317408 111486
rect 317088 111218 317130 111454
rect 317366 111218 317408 111454
rect 317088 111134 317408 111218
rect 317088 110898 317130 111134
rect 317366 110898 317408 111134
rect 317088 110866 317408 110898
rect 347808 111454 348128 111486
rect 347808 111218 347850 111454
rect 348086 111218 348128 111454
rect 347808 111134 348128 111218
rect 347808 110898 347850 111134
rect 348086 110898 348128 111134
rect 347808 110866 348128 110898
rect 378528 111454 378848 111486
rect 378528 111218 378570 111454
rect 378806 111218 378848 111454
rect 378528 111134 378848 111218
rect 378528 110898 378570 111134
rect 378806 110898 378848 111134
rect 378528 110866 378848 110898
rect 209568 93454 209888 93486
rect 209568 93218 209610 93454
rect 209846 93218 209888 93454
rect 209568 93134 209888 93218
rect 209568 92898 209610 93134
rect 209846 92898 209888 93134
rect 209568 92866 209888 92898
rect 240288 93454 240608 93486
rect 240288 93218 240330 93454
rect 240566 93218 240608 93454
rect 240288 93134 240608 93218
rect 240288 92898 240330 93134
rect 240566 92898 240608 93134
rect 240288 92866 240608 92898
rect 271008 93454 271328 93486
rect 271008 93218 271050 93454
rect 271286 93218 271328 93454
rect 271008 93134 271328 93218
rect 271008 92898 271050 93134
rect 271286 92898 271328 93134
rect 271008 92866 271328 92898
rect 301728 93454 302048 93486
rect 301728 93218 301770 93454
rect 302006 93218 302048 93454
rect 301728 93134 302048 93218
rect 301728 92898 301770 93134
rect 302006 92898 302048 93134
rect 301728 92866 302048 92898
rect 332448 93454 332768 93486
rect 332448 93218 332490 93454
rect 332726 93218 332768 93454
rect 332448 93134 332768 93218
rect 332448 92898 332490 93134
rect 332726 92898 332768 93134
rect 332448 92866 332768 92898
rect 363168 93454 363488 93486
rect 363168 93218 363210 93454
rect 363446 93218 363488 93454
rect 363168 93134 363488 93218
rect 363168 92898 363210 93134
rect 363446 92898 363488 93134
rect 363168 92866 363488 92898
rect 393888 93454 394208 93486
rect 393888 93218 393930 93454
rect 394166 93218 394208 93454
rect 393888 93134 394208 93218
rect 393888 92898 393930 93134
rect 394166 92898 394208 93134
rect 393888 92866 394208 92898
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 194208 75454 194528 75486
rect 194208 75218 194250 75454
rect 194486 75218 194528 75454
rect 194208 75134 194528 75218
rect 194208 74898 194250 75134
rect 194486 74898 194528 75134
rect 194208 74866 194528 74898
rect 224928 75454 225248 75486
rect 224928 75218 224970 75454
rect 225206 75218 225248 75454
rect 224928 75134 225248 75218
rect 224928 74898 224970 75134
rect 225206 74898 225248 75134
rect 224928 74866 225248 74898
rect 255648 75454 255968 75486
rect 255648 75218 255690 75454
rect 255926 75218 255968 75454
rect 255648 75134 255968 75218
rect 255648 74898 255690 75134
rect 255926 74898 255968 75134
rect 255648 74866 255968 74898
rect 286368 75454 286688 75486
rect 286368 75218 286410 75454
rect 286646 75218 286688 75454
rect 286368 75134 286688 75218
rect 286368 74898 286410 75134
rect 286646 74898 286688 75134
rect 286368 74866 286688 74898
rect 317088 75454 317408 75486
rect 317088 75218 317130 75454
rect 317366 75218 317408 75454
rect 317088 75134 317408 75218
rect 317088 74898 317130 75134
rect 317366 74898 317408 75134
rect 317088 74866 317408 74898
rect 347808 75454 348128 75486
rect 347808 75218 347850 75454
rect 348086 75218 348128 75454
rect 347808 75134 348128 75218
rect 347808 74898 347850 75134
rect 348086 74898 348128 75134
rect 347808 74866 348128 74898
rect 378528 75454 378848 75486
rect 378528 75218 378570 75454
rect 378806 75218 378848 75454
rect 378528 75134 378848 75218
rect 378528 74898 378570 75134
rect 378806 74898 378848 75134
rect 378528 74866 378848 74898
rect 209568 57454 209888 57486
rect 209568 57218 209610 57454
rect 209846 57218 209888 57454
rect 209568 57134 209888 57218
rect 209568 56898 209610 57134
rect 209846 56898 209888 57134
rect 209568 56866 209888 56898
rect 240288 57454 240608 57486
rect 240288 57218 240330 57454
rect 240566 57218 240608 57454
rect 240288 57134 240608 57218
rect 240288 56898 240330 57134
rect 240566 56898 240608 57134
rect 240288 56866 240608 56898
rect 271008 57454 271328 57486
rect 271008 57218 271050 57454
rect 271286 57218 271328 57454
rect 271008 57134 271328 57218
rect 271008 56898 271050 57134
rect 271286 56898 271328 57134
rect 271008 56866 271328 56898
rect 301728 57454 302048 57486
rect 301728 57218 301770 57454
rect 302006 57218 302048 57454
rect 301728 57134 302048 57218
rect 301728 56898 301770 57134
rect 302006 56898 302048 57134
rect 301728 56866 302048 56898
rect 332448 57454 332768 57486
rect 332448 57218 332490 57454
rect 332726 57218 332768 57454
rect 332448 57134 332768 57218
rect 332448 56898 332490 57134
rect 332726 56898 332768 57134
rect 332448 56866 332768 56898
rect 363168 57454 363488 57486
rect 363168 57218 363210 57454
rect 363446 57218 363488 57454
rect 363168 57134 363488 57218
rect 363168 56898 363210 57134
rect 363446 56898 363488 57134
rect 363168 56866 363488 56898
rect 393888 57454 394208 57486
rect 393888 57218 393930 57454
rect 394166 57218 394208 57454
rect 393888 57134 394208 57218
rect 393888 56898 393930 57134
rect 394166 56898 394208 57134
rect 393888 56866 394208 56898
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 194208 39454 194528 39486
rect 194208 39218 194250 39454
rect 194486 39218 194528 39454
rect 194208 39134 194528 39218
rect 194208 38898 194250 39134
rect 194486 38898 194528 39134
rect 194208 38866 194528 38898
rect 224928 39454 225248 39486
rect 224928 39218 224970 39454
rect 225206 39218 225248 39454
rect 224928 39134 225248 39218
rect 224928 38898 224970 39134
rect 225206 38898 225248 39134
rect 224928 38866 225248 38898
rect 255648 39454 255968 39486
rect 255648 39218 255690 39454
rect 255926 39218 255968 39454
rect 255648 39134 255968 39218
rect 255648 38898 255690 39134
rect 255926 38898 255968 39134
rect 255648 38866 255968 38898
rect 286368 39454 286688 39486
rect 286368 39218 286410 39454
rect 286646 39218 286688 39454
rect 286368 39134 286688 39218
rect 286368 38898 286410 39134
rect 286646 38898 286688 39134
rect 286368 38866 286688 38898
rect 317088 39454 317408 39486
rect 317088 39218 317130 39454
rect 317366 39218 317408 39454
rect 317088 39134 317408 39218
rect 317088 38898 317130 39134
rect 317366 38898 317408 39134
rect 317088 38866 317408 38898
rect 347808 39454 348128 39486
rect 347808 39218 347850 39454
rect 348086 39218 348128 39454
rect 347808 39134 348128 39218
rect 347808 38898 347850 39134
rect 348086 38898 348128 39134
rect 347808 38866 348128 38898
rect 378528 39454 378848 39486
rect 378528 39218 378570 39454
rect 378806 39218 378848 39454
rect 378528 39134 378848 39218
rect 378528 38898 378570 39134
rect 378806 38898 378848 39134
rect 378528 38866 378848 38898
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 28000
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 28000
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 28000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 28000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 28000
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 28000
rect 217794 3454 218414 28000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 7174 222134 28000
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 10894 225854 28000
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 28000
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 28000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 28000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 28000
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 28000
rect 253794 3454 254414 28000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 28000
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 28000
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 28000
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 28000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 28000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 28000
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 28000
rect 289794 3454 290414 28000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 7174 294134 28000
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 10894 297854 28000
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 28000
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 21454 308414 28000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 28000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 -5146 315854 28000
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 28000
rect 325794 3454 326414 28000
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 7174 330134 28000
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 10894 333854 28000
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 14614 337574 28000
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 21454 344414 28000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 28000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 -5146 351854 28000
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 28000
rect 361794 3454 362414 28000
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 7174 366134 28000
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 10894 369854 28000
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 14614 373574 28000
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 28000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 28000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 -5146 387854 28000
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 28000
rect 397794 3454 398414 28000
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 7174 402134 28000
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 10894 405854 28000
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 14614 409574 28000
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 132000 438134 150618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 132000 441854 154338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 132000 445574 158058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 132000 452414 164898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 132000 456134 132618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 132000 459854 136338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 132000 463574 140058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 132000 470414 146898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 132000 474134 150618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 132000 477854 154338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 132000 481574 158058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 132000 488414 164898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 132000 492134 132618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 132000 495854 136338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 132000 499574 140058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 132000 506414 146898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 132000 510134 150618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 132000 513854 154338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 132000 517574 158058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 132000 524414 164898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 132000 528134 132618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 132000 531854 136338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 132000 535574 140058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 132000 542414 146898
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 444208 111454 444528 111486
rect 444208 111218 444250 111454
rect 444486 111218 444528 111454
rect 444208 111134 444528 111218
rect 444208 110898 444250 111134
rect 444486 110898 444528 111134
rect 444208 110866 444528 110898
rect 474928 111454 475248 111486
rect 474928 111218 474970 111454
rect 475206 111218 475248 111454
rect 474928 111134 475248 111218
rect 474928 110898 474970 111134
rect 475206 110898 475248 111134
rect 474928 110866 475248 110898
rect 505648 111454 505968 111486
rect 505648 111218 505690 111454
rect 505926 111218 505968 111454
rect 505648 111134 505968 111218
rect 505648 110898 505690 111134
rect 505926 110898 505968 111134
rect 505648 110866 505968 110898
rect 536368 111454 536688 111486
rect 536368 111218 536410 111454
rect 536646 111218 536688 111454
rect 536368 111134 536688 111218
rect 536368 110898 536410 111134
rect 536646 110898 536688 111134
rect 536368 110866 536688 110898
rect 459568 93454 459888 93486
rect 459568 93218 459610 93454
rect 459846 93218 459888 93454
rect 459568 93134 459888 93218
rect 459568 92898 459610 93134
rect 459846 92898 459888 93134
rect 459568 92866 459888 92898
rect 490288 93454 490608 93486
rect 490288 93218 490330 93454
rect 490566 93218 490608 93454
rect 490288 93134 490608 93218
rect 490288 92898 490330 93134
rect 490566 92898 490608 93134
rect 490288 92866 490608 92898
rect 521008 93454 521328 93486
rect 521008 93218 521050 93454
rect 521286 93218 521328 93454
rect 521008 93134 521328 93218
rect 521008 92898 521050 93134
rect 521286 92898 521328 93134
rect 521008 92866 521328 92898
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 444208 75454 444528 75486
rect 444208 75218 444250 75454
rect 444486 75218 444528 75454
rect 444208 75134 444528 75218
rect 444208 74898 444250 75134
rect 444486 74898 444528 75134
rect 444208 74866 444528 74898
rect 474928 75454 475248 75486
rect 474928 75218 474970 75454
rect 475206 75218 475248 75454
rect 474928 75134 475248 75218
rect 474928 74898 474970 75134
rect 475206 74898 475248 75134
rect 474928 74866 475248 74898
rect 505648 75454 505968 75486
rect 505648 75218 505690 75454
rect 505926 75218 505968 75454
rect 505648 75134 505968 75218
rect 505648 74898 505690 75134
rect 505926 74898 505968 75134
rect 505648 74866 505968 74898
rect 536368 75454 536688 75486
rect 536368 75218 536410 75454
rect 536646 75218 536688 75454
rect 536368 75134 536688 75218
rect 536368 74898 536410 75134
rect 536646 74898 536688 75134
rect 536368 74866 536688 74898
rect 459568 57454 459888 57486
rect 459568 57218 459610 57454
rect 459846 57218 459888 57454
rect 459568 57134 459888 57218
rect 459568 56898 459610 57134
rect 459846 56898 459888 57134
rect 459568 56866 459888 56898
rect 490288 57454 490608 57486
rect 490288 57218 490330 57454
rect 490566 57218 490608 57454
rect 490288 57134 490608 57218
rect 490288 56898 490330 57134
rect 490566 56898 490608 57134
rect 490288 56866 490608 56898
rect 521008 57454 521328 57486
rect 521008 57218 521050 57454
rect 521286 57218 521328 57454
rect 521008 57134 521328 57218
rect 521008 56898 521050 57134
rect 521286 56898 521328 57134
rect 521008 56866 521328 56898
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 444208 39454 444528 39486
rect 444208 39218 444250 39454
rect 444486 39218 444528 39454
rect 444208 39134 444528 39218
rect 444208 38898 444250 39134
rect 444486 38898 444528 39134
rect 444208 38866 444528 38898
rect 474928 39454 475248 39486
rect 474928 39218 474970 39454
rect 475206 39218 475248 39454
rect 474928 39134 475248 39218
rect 474928 38898 474970 39134
rect 475206 38898 475248 39134
rect 474928 38866 475248 38898
rect 505648 39454 505968 39486
rect 505648 39218 505690 39454
rect 505926 39218 505968 39454
rect 505648 39134 505968 39218
rect 505648 38898 505690 39134
rect 505926 38898 505968 39134
rect 505648 38866 505968 38898
rect 536368 39454 536688 39486
rect 536368 39218 536410 39454
rect 536646 39218 536688 39454
rect 536368 39134 536688 39218
rect 536368 38898 536410 39134
rect 536646 38898 536688 39134
rect 536368 38866 536688 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 7174 438134 28000
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 10894 441854 28000
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 14614 445574 28000
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 21454 452414 28000
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 28000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 -5146 459854 28000
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 28000
rect 469794 3454 470414 28000
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 7174 474134 28000
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 10894 477854 28000
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 14614 481574 28000
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 21454 488414 28000
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 28000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 -5146 495854 28000
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 28000
rect 505794 3454 506414 28000
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 7174 510134 28000
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 10894 513854 28000
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 14614 517574 28000
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 21454 524414 28000
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 25174 528134 28000
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 -5146 531854 28000
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 28000
rect 541794 3454 542414 28000
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 51008 363218 51244 363454
rect 51008 362898 51244 363134
rect 144712 363218 144948 363454
rect 144712 362898 144948 363134
rect 50328 345218 50564 345454
rect 50328 344898 50564 345134
rect 145392 345218 145628 345454
rect 145392 344898 145628 345134
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 51008 327218 51244 327454
rect 51008 326898 51244 327134
rect 144712 327218 144948 327454
rect 144712 326898 144948 327134
rect 50328 309218 50564 309454
rect 50328 308898 50564 309134
rect 145392 309218 145628 309454
rect 145392 308898 145628 309134
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 34250 111218 34486 111454
rect 34250 110898 34486 111134
rect 64970 111218 65206 111454
rect 64970 110898 65206 111134
rect 95690 111218 95926 111454
rect 95690 110898 95926 111134
rect 126410 111218 126646 111454
rect 126410 110898 126646 111134
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 49610 93218 49846 93454
rect 49610 92898 49846 93134
rect 80330 93218 80566 93454
rect 80330 92898 80566 93134
rect 111050 93218 111286 93454
rect 111050 92898 111286 93134
rect 34250 75218 34486 75454
rect 34250 74898 34486 75134
rect 64970 75218 65206 75454
rect 64970 74898 65206 75134
rect 95690 75218 95926 75454
rect 95690 74898 95926 75134
rect 126410 75218 126646 75454
rect 126410 74898 126646 75134
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 49610 57218 49846 57454
rect 49610 56898 49846 57134
rect 80330 57218 80566 57454
rect 80330 56898 80566 57134
rect 111050 57218 111286 57454
rect 111050 56898 111286 57134
rect 34250 39218 34486 39454
rect 34250 38898 34486 39134
rect 64970 39218 65206 39454
rect 64970 38898 65206 39134
rect 95690 39218 95926 39454
rect 95690 38898 95926 39134
rect 126410 39218 126646 39454
rect 126410 38898 126646 39134
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 211008 363218 211244 363454
rect 211008 362898 211244 363134
rect 304712 363218 304948 363454
rect 304712 362898 304948 363134
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 210328 345218 210564 345454
rect 210328 344898 210564 345134
rect 305392 345218 305628 345454
rect 305392 344898 305628 345134
rect 211008 327218 211244 327454
rect 211008 326898 211244 327134
rect 304712 327218 304948 327454
rect 304712 326898 304948 327134
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 210328 309218 210564 309454
rect 210328 308898 210564 309134
rect 305392 309218 305628 309454
rect 305392 308898 305628 309134
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 209610 237218 209846 237454
rect 209610 236898 209846 237134
rect 240330 237218 240566 237454
rect 240330 236898 240566 237134
rect 271050 237218 271286 237454
rect 271050 236898 271286 237134
rect 301770 237218 302006 237454
rect 301770 236898 302006 237134
rect 332490 237218 332726 237454
rect 332490 236898 332726 237134
rect 363210 237218 363446 237454
rect 363210 236898 363446 237134
rect 393930 237218 394166 237454
rect 393930 236898 394166 237134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 194250 219218 194486 219454
rect 194250 218898 194486 219134
rect 224970 219218 225206 219454
rect 224970 218898 225206 219134
rect 255690 219218 255926 219454
rect 255690 218898 255926 219134
rect 286410 219218 286646 219454
rect 286410 218898 286646 219134
rect 317130 219218 317366 219454
rect 317130 218898 317366 219134
rect 347850 219218 348086 219454
rect 347850 218898 348086 219134
rect 378570 219218 378806 219454
rect 378570 218898 378806 219134
rect 209610 201218 209846 201454
rect 209610 200898 209846 201134
rect 240330 201218 240566 201454
rect 240330 200898 240566 201134
rect 271050 201218 271286 201454
rect 271050 200898 271286 201134
rect 301770 201218 302006 201454
rect 301770 200898 302006 201134
rect 332490 201218 332726 201454
rect 332490 200898 332726 201134
rect 363210 201218 363446 201454
rect 363210 200898 363446 201134
rect 393930 201218 394166 201454
rect 393930 200898 394166 201134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 194250 183218 194486 183454
rect 194250 182898 194486 183134
rect 224970 183218 225206 183454
rect 224970 182898 225206 183134
rect 255690 183218 255926 183454
rect 255690 182898 255926 183134
rect 286410 183218 286646 183454
rect 286410 182898 286646 183134
rect 317130 183218 317366 183454
rect 317130 182898 317366 183134
rect 347850 183218 348086 183454
rect 347850 182898 348086 183134
rect 378570 183218 378806 183454
rect 378570 182898 378806 183134
rect 209610 165218 209846 165454
rect 209610 164898 209846 165134
rect 240330 165218 240566 165454
rect 240330 164898 240566 165134
rect 271050 165218 271286 165454
rect 271050 164898 271286 165134
rect 301770 165218 302006 165454
rect 301770 164898 302006 165134
rect 332490 165218 332726 165454
rect 332490 164898 332726 165134
rect 363210 165218 363446 165454
rect 363210 164898 363446 165134
rect 393930 165218 394166 165454
rect 393930 164898 394166 165134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 194250 147218 194486 147454
rect 194250 146898 194486 147134
rect 224970 147218 225206 147454
rect 224970 146898 225206 147134
rect 255690 147218 255926 147454
rect 255690 146898 255926 147134
rect 286410 147218 286646 147454
rect 286410 146898 286646 147134
rect 317130 147218 317366 147454
rect 317130 146898 317366 147134
rect 347850 147218 348086 147454
rect 347850 146898 348086 147134
rect 378570 147218 378806 147454
rect 378570 146898 378806 147134
rect 209610 129218 209846 129454
rect 209610 128898 209846 129134
rect 240330 129218 240566 129454
rect 240330 128898 240566 129134
rect 271050 129218 271286 129454
rect 271050 128898 271286 129134
rect 301770 129218 302006 129454
rect 301770 128898 302006 129134
rect 332490 129218 332726 129454
rect 332490 128898 332726 129134
rect 363210 129218 363446 129454
rect 363210 128898 363446 129134
rect 393930 129218 394166 129454
rect 393930 128898 394166 129134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 194250 111218 194486 111454
rect 194250 110898 194486 111134
rect 224970 111218 225206 111454
rect 224970 110898 225206 111134
rect 255690 111218 255926 111454
rect 255690 110898 255926 111134
rect 286410 111218 286646 111454
rect 286410 110898 286646 111134
rect 317130 111218 317366 111454
rect 317130 110898 317366 111134
rect 347850 111218 348086 111454
rect 347850 110898 348086 111134
rect 378570 111218 378806 111454
rect 378570 110898 378806 111134
rect 209610 93218 209846 93454
rect 209610 92898 209846 93134
rect 240330 93218 240566 93454
rect 240330 92898 240566 93134
rect 271050 93218 271286 93454
rect 271050 92898 271286 93134
rect 301770 93218 302006 93454
rect 301770 92898 302006 93134
rect 332490 93218 332726 93454
rect 332490 92898 332726 93134
rect 363210 93218 363446 93454
rect 363210 92898 363446 93134
rect 393930 93218 394166 93454
rect 393930 92898 394166 93134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 194250 75218 194486 75454
rect 194250 74898 194486 75134
rect 224970 75218 225206 75454
rect 224970 74898 225206 75134
rect 255690 75218 255926 75454
rect 255690 74898 255926 75134
rect 286410 75218 286646 75454
rect 286410 74898 286646 75134
rect 317130 75218 317366 75454
rect 317130 74898 317366 75134
rect 347850 75218 348086 75454
rect 347850 74898 348086 75134
rect 378570 75218 378806 75454
rect 378570 74898 378806 75134
rect 209610 57218 209846 57454
rect 209610 56898 209846 57134
rect 240330 57218 240566 57454
rect 240330 56898 240566 57134
rect 271050 57218 271286 57454
rect 271050 56898 271286 57134
rect 301770 57218 302006 57454
rect 301770 56898 302006 57134
rect 332490 57218 332726 57454
rect 332490 56898 332726 57134
rect 363210 57218 363446 57454
rect 363210 56898 363446 57134
rect 393930 57218 394166 57454
rect 393930 56898 394166 57134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 194250 39218 194486 39454
rect 194250 38898 194486 39134
rect 224970 39218 225206 39454
rect 224970 38898 225206 39134
rect 255690 39218 255926 39454
rect 255690 38898 255926 39134
rect 286410 39218 286646 39454
rect 286410 38898 286646 39134
rect 317130 39218 317366 39454
rect 317130 38898 317366 39134
rect 347850 39218 348086 39454
rect 347850 38898 348086 39134
rect 378570 39218 378806 39454
rect 378570 38898 378806 39134
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 444250 111218 444486 111454
rect 444250 110898 444486 111134
rect 474970 111218 475206 111454
rect 474970 110898 475206 111134
rect 505690 111218 505926 111454
rect 505690 110898 505926 111134
rect 536410 111218 536646 111454
rect 536410 110898 536646 111134
rect 459610 93218 459846 93454
rect 459610 92898 459846 93134
rect 490330 93218 490566 93454
rect 490330 92898 490566 93134
rect 521050 93218 521286 93454
rect 521050 92898 521286 93134
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 444250 75218 444486 75454
rect 444250 74898 444486 75134
rect 474970 75218 475206 75454
rect 474970 74898 475206 75134
rect 505690 75218 505926 75454
rect 505690 74898 505926 75134
rect 536410 75218 536646 75454
rect 536410 74898 536646 75134
rect 459610 57218 459846 57454
rect 459610 56898 459846 57134
rect 490330 57218 490566 57454
rect 490330 56898 490566 57134
rect 521050 57218 521286 57454
rect 521050 56898 521286 57134
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 444250 39218 444486 39454
rect 444250 38898 444486 39134
rect 474970 39218 475206 39454
rect 474970 38898 475206 39134
rect 505690 39218 505926 39454
rect 505690 38898 505926 39134
rect 536410 39218 536646 39454
rect 536410 38898 536646 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 51008 363454
rect 51244 363218 144712 363454
rect 144948 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 211008 363454
rect 211244 363218 304712 363454
rect 304948 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 51008 363134
rect 51244 362898 144712 363134
rect 144948 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 211008 363134
rect 211244 362898 304712 363134
rect 304948 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 50328 345454
rect 50564 345218 145392 345454
rect 145628 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 210328 345454
rect 210564 345218 305392 345454
rect 305628 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 50328 345134
rect 50564 344898 145392 345134
rect 145628 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 210328 345134
rect 210564 344898 305392 345134
rect 305628 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 51008 327454
rect 51244 327218 144712 327454
rect 144948 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 211008 327454
rect 211244 327218 304712 327454
rect 304948 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 51008 327134
rect 51244 326898 144712 327134
rect 144948 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 211008 327134
rect 211244 326898 304712 327134
rect 304948 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 50328 309454
rect 50564 309218 145392 309454
rect 145628 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 210328 309454
rect 210564 309218 305392 309454
rect 305628 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 50328 309134
rect 50564 308898 145392 309134
rect 145628 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 210328 309134
rect 210564 308898 305392 309134
rect 305628 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 209610 237454
rect 209846 237218 240330 237454
rect 240566 237218 271050 237454
rect 271286 237218 301770 237454
rect 302006 237218 332490 237454
rect 332726 237218 363210 237454
rect 363446 237218 393930 237454
rect 394166 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 209610 237134
rect 209846 236898 240330 237134
rect 240566 236898 271050 237134
rect 271286 236898 301770 237134
rect 302006 236898 332490 237134
rect 332726 236898 363210 237134
rect 363446 236898 393930 237134
rect 394166 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 194250 219454
rect 194486 219218 224970 219454
rect 225206 219218 255690 219454
rect 255926 219218 286410 219454
rect 286646 219218 317130 219454
rect 317366 219218 347850 219454
rect 348086 219218 378570 219454
rect 378806 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 194250 219134
rect 194486 218898 224970 219134
rect 225206 218898 255690 219134
rect 255926 218898 286410 219134
rect 286646 218898 317130 219134
rect 317366 218898 347850 219134
rect 348086 218898 378570 219134
rect 378806 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 209610 201454
rect 209846 201218 240330 201454
rect 240566 201218 271050 201454
rect 271286 201218 301770 201454
rect 302006 201218 332490 201454
rect 332726 201218 363210 201454
rect 363446 201218 393930 201454
rect 394166 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 209610 201134
rect 209846 200898 240330 201134
rect 240566 200898 271050 201134
rect 271286 200898 301770 201134
rect 302006 200898 332490 201134
rect 332726 200898 363210 201134
rect 363446 200898 393930 201134
rect 394166 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 194250 183454
rect 194486 183218 224970 183454
rect 225206 183218 255690 183454
rect 255926 183218 286410 183454
rect 286646 183218 317130 183454
rect 317366 183218 347850 183454
rect 348086 183218 378570 183454
rect 378806 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 194250 183134
rect 194486 182898 224970 183134
rect 225206 182898 255690 183134
rect 255926 182898 286410 183134
rect 286646 182898 317130 183134
rect 317366 182898 347850 183134
rect 348086 182898 378570 183134
rect 378806 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 209610 165454
rect 209846 165218 240330 165454
rect 240566 165218 271050 165454
rect 271286 165218 301770 165454
rect 302006 165218 332490 165454
rect 332726 165218 363210 165454
rect 363446 165218 393930 165454
rect 394166 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 209610 165134
rect 209846 164898 240330 165134
rect 240566 164898 271050 165134
rect 271286 164898 301770 165134
rect 302006 164898 332490 165134
rect 332726 164898 363210 165134
rect 363446 164898 393930 165134
rect 394166 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 194250 147454
rect 194486 147218 224970 147454
rect 225206 147218 255690 147454
rect 255926 147218 286410 147454
rect 286646 147218 317130 147454
rect 317366 147218 347850 147454
rect 348086 147218 378570 147454
rect 378806 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 194250 147134
rect 194486 146898 224970 147134
rect 225206 146898 255690 147134
rect 255926 146898 286410 147134
rect 286646 146898 317130 147134
rect 317366 146898 347850 147134
rect 348086 146898 378570 147134
rect 378806 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 209610 129454
rect 209846 129218 240330 129454
rect 240566 129218 271050 129454
rect 271286 129218 301770 129454
rect 302006 129218 332490 129454
rect 332726 129218 363210 129454
rect 363446 129218 393930 129454
rect 394166 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 209610 129134
rect 209846 128898 240330 129134
rect 240566 128898 271050 129134
rect 271286 128898 301770 129134
rect 302006 128898 332490 129134
rect 332726 128898 363210 129134
rect 363446 128898 393930 129134
rect 394166 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 34250 111454
rect 34486 111218 64970 111454
rect 65206 111218 95690 111454
rect 95926 111218 126410 111454
rect 126646 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 194250 111454
rect 194486 111218 224970 111454
rect 225206 111218 255690 111454
rect 255926 111218 286410 111454
rect 286646 111218 317130 111454
rect 317366 111218 347850 111454
rect 348086 111218 378570 111454
rect 378806 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 444250 111454
rect 444486 111218 474970 111454
rect 475206 111218 505690 111454
rect 505926 111218 536410 111454
rect 536646 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 34250 111134
rect 34486 110898 64970 111134
rect 65206 110898 95690 111134
rect 95926 110898 126410 111134
rect 126646 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 194250 111134
rect 194486 110898 224970 111134
rect 225206 110898 255690 111134
rect 255926 110898 286410 111134
rect 286646 110898 317130 111134
rect 317366 110898 347850 111134
rect 348086 110898 378570 111134
rect 378806 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 444250 111134
rect 444486 110898 474970 111134
rect 475206 110898 505690 111134
rect 505926 110898 536410 111134
rect 536646 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 49610 93454
rect 49846 93218 80330 93454
rect 80566 93218 111050 93454
rect 111286 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 209610 93454
rect 209846 93218 240330 93454
rect 240566 93218 271050 93454
rect 271286 93218 301770 93454
rect 302006 93218 332490 93454
rect 332726 93218 363210 93454
rect 363446 93218 393930 93454
rect 394166 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 459610 93454
rect 459846 93218 490330 93454
rect 490566 93218 521050 93454
rect 521286 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 49610 93134
rect 49846 92898 80330 93134
rect 80566 92898 111050 93134
rect 111286 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 209610 93134
rect 209846 92898 240330 93134
rect 240566 92898 271050 93134
rect 271286 92898 301770 93134
rect 302006 92898 332490 93134
rect 332726 92898 363210 93134
rect 363446 92898 393930 93134
rect 394166 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 459610 93134
rect 459846 92898 490330 93134
rect 490566 92898 521050 93134
rect 521286 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 34250 75454
rect 34486 75218 64970 75454
rect 65206 75218 95690 75454
rect 95926 75218 126410 75454
rect 126646 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 194250 75454
rect 194486 75218 224970 75454
rect 225206 75218 255690 75454
rect 255926 75218 286410 75454
rect 286646 75218 317130 75454
rect 317366 75218 347850 75454
rect 348086 75218 378570 75454
rect 378806 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 444250 75454
rect 444486 75218 474970 75454
rect 475206 75218 505690 75454
rect 505926 75218 536410 75454
rect 536646 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 34250 75134
rect 34486 74898 64970 75134
rect 65206 74898 95690 75134
rect 95926 74898 126410 75134
rect 126646 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 194250 75134
rect 194486 74898 224970 75134
rect 225206 74898 255690 75134
rect 255926 74898 286410 75134
rect 286646 74898 317130 75134
rect 317366 74898 347850 75134
rect 348086 74898 378570 75134
rect 378806 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 444250 75134
rect 444486 74898 474970 75134
rect 475206 74898 505690 75134
rect 505926 74898 536410 75134
rect 536646 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 49610 57454
rect 49846 57218 80330 57454
rect 80566 57218 111050 57454
rect 111286 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 209610 57454
rect 209846 57218 240330 57454
rect 240566 57218 271050 57454
rect 271286 57218 301770 57454
rect 302006 57218 332490 57454
rect 332726 57218 363210 57454
rect 363446 57218 393930 57454
rect 394166 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 459610 57454
rect 459846 57218 490330 57454
rect 490566 57218 521050 57454
rect 521286 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 49610 57134
rect 49846 56898 80330 57134
rect 80566 56898 111050 57134
rect 111286 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 209610 57134
rect 209846 56898 240330 57134
rect 240566 56898 271050 57134
rect 271286 56898 301770 57134
rect 302006 56898 332490 57134
rect 332726 56898 363210 57134
rect 363446 56898 393930 57134
rect 394166 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 459610 57134
rect 459846 56898 490330 57134
rect 490566 56898 521050 57134
rect 521286 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 34250 39454
rect 34486 39218 64970 39454
rect 65206 39218 95690 39454
rect 95926 39218 126410 39454
rect 126646 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 194250 39454
rect 194486 39218 224970 39454
rect 225206 39218 255690 39454
rect 255926 39218 286410 39454
rect 286646 39218 317130 39454
rect 317366 39218 347850 39454
rect 348086 39218 378570 39454
rect 378806 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 444250 39454
rect 444486 39218 474970 39454
rect 475206 39218 505690 39454
rect 505926 39218 536410 39454
rect 536646 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 34250 39134
rect 34486 38898 64970 39134
rect 65206 38898 95690 39134
rect 95926 38898 126410 39134
rect 126646 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 194250 39134
rect 194486 38898 224970 39134
rect 225206 38898 255690 39134
rect 255926 38898 286410 39134
rect 286646 38898 317130 39134
rect 317366 38898 347850 39134
rect 348086 38898 378570 39134
rect 378806 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 444250 39134
rect 444486 38898 474970 39134
rect 475206 38898 505690 39134
rect 505926 38898 536410 39134
rect 536646 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use Core  core
timestamp 0
transform 1 0 30000 0 1 30000
box 1066 0 100000 100000
use sky130_sram_1kbyte_1rw1r_32x256_8  dmem
timestamp 0
transform 1 0 210000 0 1 300000
box 0 0 95956 79500
use sky130_sram_1kbyte_1rw1r_32x256_8  imem
timestamp 0
transform 1 0 50000 0 1 300000
box 0 0 95956 79500
use Motor_Top  motor
timestamp 0
transform 1 0 440000 0 1 30000
box 0 0 100000 100000
use WB_InterConnect  wb_inter_connect
timestamp 0
transform 1 0 190000 0 1 30000
box 0 0 220000 220000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 132000 74414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 132000 110414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 252000 218414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 252000 254414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 252000 290414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 132000 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 381500 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 381500 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 381500 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 381500 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 381500 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 381500 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 252000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 252000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 252000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 132000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 132000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 132000 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 132000 78134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 132000 114134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 252000 222134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 252000 258134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 252000 294134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 132000 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 381500 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 381500 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 381500 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 381500 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 381500 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 252000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 252000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 252000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 132000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 132000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 132000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 132000 81854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 132000 117854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 252000 225854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 252000 261854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 252000 297854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 132000 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 381500 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 381500 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 252000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 381500 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 381500 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 381500 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 252000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 252000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 252000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 132000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 132000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 132000 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 132000 49574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 132000 85574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 132000 121574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 252000 229574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 252000 265574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 252000 301574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 381500 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 381500 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 381500 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 252000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 381500 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 381500 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 381500 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 252000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 252000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 252000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 132000 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 132000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 132000 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 132000 63854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 132000 99854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 252000 243854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 252000 279854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 381500 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 381500 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 381500 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 252000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 381500 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 381500 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 252000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 252000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 252000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 132000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 132000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 132000 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 132000 67574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 132000 103574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 252000 211574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 252000 247574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 252000 283574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 132000 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 381500 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 381500 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 381500 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 381500 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 381500 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 381500 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 252000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 252000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 252000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 132000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 132000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 132000 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 132000 56414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 132000 92414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 132000 128414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 252000 236414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 252000 272414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 252000 308414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 381500 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 381500 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 381500 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 252000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 381500 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 381500 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 381500 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 252000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 252000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 132000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 132000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 132000 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 132000 60134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 132000 96134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 132000 132134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 252000 240134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 252000 276134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 381500 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 381500 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 381500 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 252000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 381500 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 381500 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 252000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 252000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 252000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 132000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 132000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 132000 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
