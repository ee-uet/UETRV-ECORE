VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Motor_Top
  CLASS BLOCK ;
  FOREIGN Motor_Top ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END clock
  PIN io_ba_match
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 496.000 41.770 500.000 ;
    END
  END io_ba_match
  PIN io_motor_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END io_motor_irq
  PIN io_pwm_high
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 496.000 8.650 500.000 ;
    END
  END io_pwm_high
  PIN io_pwm_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 496.000 25.210 500.000 ;
    END
  END io_pwm_low
  PIN io_qei_ch_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 8.200 500.000 8.800 ;
    END
  END io_qei_ch_a
  PIN io_qei_ch_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 496.000 58.330 500.000 ;
    END
  END io_qei_ch_b
  PIN io_wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 25.200 500.000 25.800 ;
    END
  END io_wbs_ack_o
  PIN io_wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 76.880 500.000 77.480 ;
    END
  END io_wbs_data_o[0]
  PIN io_wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END io_wbs_data_o[10]
  PIN io_wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END io_wbs_data_o[11]
  PIN io_wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 496.000 274.990 500.000 ;
    END
  END io_wbs_data_o[12]
  PIN io_wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END io_wbs_data_o[13]
  PIN io_wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 496.000 291.550 500.000 ;
    END
  END io_wbs_data_o[14]
  PIN io_wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END io_wbs_data_o[15]
  PIN io_wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END io_wbs_data_o[16]
  PIN io_wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 335.280 500.000 335.880 ;
    END
  END io_wbs_data_o[17]
  PIN io_wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END io_wbs_data_o[18]
  PIN io_wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END io_wbs_data_o[19]
  PIN io_wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END io_wbs_data_o[1]
  PIN io_wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END io_wbs_data_o[20]
  PIN io_wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 496.000 391.830 500.000 ;
    END
  END io_wbs_data_o[21]
  PIN io_wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END io_wbs_data_o[22]
  PIN io_wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END io_wbs_data_o[23]
  PIN io_wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 4.000 ;
    END
  END io_wbs_data_o[24]
  PIN io_wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 496.000 441.970 500.000 ;
    END
  END io_wbs_data_o[25]
  PIN io_wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 421.640 500.000 422.240 ;
    END
  END io_wbs_data_o[26]
  PIN io_wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 496.000 458.530 500.000 ;
    END
  END io_wbs_data_o[27]
  PIN io_wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 496.000 475.090 500.000 ;
    END
  END io_wbs_data_o[28]
  PIN io_wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END io_wbs_data_o[29]
  PIN io_wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 496.000 91.910 500.000 ;
    END
  END io_wbs_data_o[2]
  PIN io_wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END io_wbs_data_o[30]
  PIN io_wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 473.320 500.000 473.920 ;
    END
  END io_wbs_data_o[31]
  PIN io_wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 496.000 108.470 500.000 ;
    END
  END io_wbs_data_o[3]
  PIN io_wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 496.000 141.590 500.000 ;
    END
  END io_wbs_data_o[4]
  PIN io_wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.960 4.000 183.560 ;
    END
  END io_wbs_data_o[5]
  PIN io_wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 163.240 500.000 163.840 ;
    END
  END io_wbs_data_o[6]
  PIN io_wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 496.000 191.730 500.000 ;
    END
  END io_wbs_data_o[7]
  PIN io_wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END io_wbs_data_o[8]
  PIN io_wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 231.920 500.000 232.520 ;
    END
  END io_wbs_data_o[9]
  PIN io_wbs_m2s_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END io_wbs_m2s_addr[0]
  PIN io_wbs_m2s_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END io_wbs_m2s_addr[10]
  PIN io_wbs_m2s_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 266.600 500.000 267.200 ;
    END
  END io_wbs_m2s_addr[11]
  PIN io_wbs_m2s_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END io_wbs_m2s_addr[12]
  PIN io_wbs_m2s_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 283.600 500.000 284.200 ;
    END
  END io_wbs_m2s_addr[13]
  PIN io_wbs_m2s_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 496.000 308.570 500.000 ;
    END
  END io_wbs_m2s_addr[14]
  PIN io_wbs_m2s_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 496.000 341.690 500.000 ;
    END
  END io_wbs_m2s_addr[15]
  PIN io_wbs_m2s_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 93.880 500.000 94.480 ;
    END
  END io_wbs_m2s_addr[1]
  PIN io_wbs_m2s_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END io_wbs_m2s_addr[2]
  PIN io_wbs_m2s_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 496.000 125.030 500.000 ;
    END
  END io_wbs_m2s_addr[3]
  PIN io_wbs_m2s_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 496.000 158.610 500.000 ;
    END
  END io_wbs_m2s_addr[4]
  PIN io_wbs_m2s_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 145.560 500.000 146.160 ;
    END
  END io_wbs_m2s_addr[5]
  PIN io_wbs_m2s_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 180.240 500.000 180.840 ;
    END
  END io_wbs_m2s_addr[6]
  PIN io_wbs_m2s_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 496.000 208.290 500.000 ;
    END
  END io_wbs_m2s_addr[7]
  PIN io_wbs_m2s_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 496.000 225.310 500.000 ;
    END
  END io_wbs_m2s_addr[8]
  PIN io_wbs_m2s_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 248.920 500.000 249.520 ;
    END
  END io_wbs_m2s_addr[9]
  PIN io_wbs_m2s_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 496.000 74.890 500.000 ;
    END
  END io_wbs_m2s_data[0]
  PIN io_wbs_m2s_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END io_wbs_m2s_data[10]
  PIN io_wbs_m2s_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 496.000 258.430 500.000 ;
    END
  END io_wbs_m2s_data[11]
  PIN io_wbs_m2s_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END io_wbs_m2s_data[12]
  PIN io_wbs_m2s_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 300.600 500.000 301.200 ;
    END
  END io_wbs_m2s_data[13]
  PIN io_wbs_m2s_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 496.000 325.130 500.000 ;
    END
  END io_wbs_m2s_data[14]
  PIN io_wbs_m2s_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 318.280 500.000 318.880 ;
    END
  END io_wbs_m2s_data[15]
  PIN io_wbs_m2s_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 496.000 358.250 500.000 ;
    END
  END io_wbs_m2s_data[16]
  PIN io_wbs_m2s_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 496.000 375.270 500.000 ;
    END
  END io_wbs_m2s_data[17]
  PIN io_wbs_m2s_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 352.280 500.000 352.880 ;
    END
  END io_wbs_m2s_data[18]
  PIN io_wbs_m2s_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 369.960 500.000 370.560 ;
    END
  END io_wbs_m2s_data[19]
  PIN io_wbs_m2s_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END io_wbs_m2s_data[1]
  PIN io_wbs_m2s_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END io_wbs_m2s_data[20]
  PIN io_wbs_m2s_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 386.960 500.000 387.560 ;
    END
  END io_wbs_m2s_data[21]
  PIN io_wbs_m2s_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 496.000 408.390 500.000 ;
    END
  END io_wbs_m2s_data[22]
  PIN io_wbs_m2s_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 496.000 424.950 500.000 ;
    END
  END io_wbs_m2s_data[23]
  PIN io_wbs_m2s_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END io_wbs_m2s_data[24]
  PIN io_wbs_m2s_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 403.960 500.000 404.560 ;
    END
  END io_wbs_m2s_data[25]
  PIN io_wbs_m2s_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END io_wbs_m2s_data[26]
  PIN io_wbs_m2s_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 438.640 500.000 439.240 ;
    END
  END io_wbs_m2s_data[27]
  PIN io_wbs_m2s_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 455.640 500.000 456.240 ;
    END
  END io_wbs_m2s_data[28]
  PIN io_wbs_m2s_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END io_wbs_m2s_data[29]
  PIN io_wbs_m2s_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 128.560 500.000 129.160 ;
    END
  END io_wbs_m2s_data[2]
  PIN io_wbs_m2s_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 496.000 491.650 500.000 ;
    END
  END io_wbs_m2s_data[30]
  PIN io_wbs_m2s_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 490.320 500.000 490.920 ;
    END
  END io_wbs_m2s_data[31]
  PIN io_wbs_m2s_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END io_wbs_m2s_data[3]
  PIN io_wbs_m2s_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 496.000 175.170 500.000 ;
    END
  END io_wbs_m2s_data[4]
  PIN io_wbs_m2s_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END io_wbs_m2s_data[5]
  PIN io_wbs_m2s_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END io_wbs_m2s_data[6]
  PIN io_wbs_m2s_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 197.240 500.000 197.840 ;
    END
  END io_wbs_m2s_data[7]
  PIN io_wbs_m2s_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 214.920 500.000 215.520 ;
    END
  END io_wbs_m2s_data[8]
  PIN io_wbs_m2s_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 496.000 241.870 500.000 ;
    END
  END io_wbs_m2s_data[9]
  PIN io_wbs_m2s_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END io_wbs_m2s_sel[0]
  PIN io_wbs_m2s_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 111.560 500.000 112.160 ;
    END
  END io_wbs_m2s_sel[1]
  PIN io_wbs_m2s_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END io_wbs_m2s_sel[2]
  PIN io_wbs_m2s_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END io_wbs_m2s_sel[3]
  PIN io_wbs_m2s_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 42.200 500.000 42.800 ;
    END
  END io_wbs_m2s_stb
  PIN io_wbs_m2s_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 59.880 500.000 60.480 ;
    END
  END io_wbs_m2s_we
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 5.520 10.240 494.040 487.120 ;
      LAYER met2 ;
        RECT 6.990 495.720 8.090 496.810 ;
        RECT 8.930 495.720 24.650 496.810 ;
        RECT 25.490 495.720 41.210 496.810 ;
        RECT 42.050 495.720 57.770 496.810 ;
        RECT 58.610 495.720 74.330 496.810 ;
        RECT 75.170 495.720 91.350 496.810 ;
        RECT 92.190 495.720 107.910 496.810 ;
        RECT 108.750 495.720 124.470 496.810 ;
        RECT 125.310 495.720 141.030 496.810 ;
        RECT 141.870 495.720 158.050 496.810 ;
        RECT 158.890 495.720 174.610 496.810 ;
        RECT 175.450 495.720 191.170 496.810 ;
        RECT 192.010 495.720 207.730 496.810 ;
        RECT 208.570 495.720 224.750 496.810 ;
        RECT 225.590 495.720 241.310 496.810 ;
        RECT 242.150 495.720 257.870 496.810 ;
        RECT 258.710 495.720 274.430 496.810 ;
        RECT 275.270 495.720 290.990 496.810 ;
        RECT 291.830 495.720 308.010 496.810 ;
        RECT 308.850 495.720 324.570 496.810 ;
        RECT 325.410 495.720 341.130 496.810 ;
        RECT 341.970 495.720 357.690 496.810 ;
        RECT 358.530 495.720 374.710 496.810 ;
        RECT 375.550 495.720 391.270 496.810 ;
        RECT 392.110 495.720 407.830 496.810 ;
        RECT 408.670 495.720 424.390 496.810 ;
        RECT 425.230 495.720 441.410 496.810 ;
        RECT 442.250 495.720 457.970 496.810 ;
        RECT 458.810 495.720 474.530 496.810 ;
        RECT 475.370 495.720 491.090 496.810 ;
        RECT 6.990 4.280 491.650 495.720 ;
        RECT 6.990 3.670 11.310 4.280 ;
        RECT 12.150 3.670 34.770 4.280 ;
        RECT 35.610 3.670 58.690 4.280 ;
        RECT 59.530 3.670 82.610 4.280 ;
        RECT 83.450 3.670 106.530 4.280 ;
        RECT 107.370 3.670 129.990 4.280 ;
        RECT 130.830 3.670 153.910 4.280 ;
        RECT 154.750 3.670 177.830 4.280 ;
        RECT 178.670 3.670 201.750 4.280 ;
        RECT 202.590 3.670 225.210 4.280 ;
        RECT 226.050 3.670 249.130 4.280 ;
        RECT 249.970 3.670 273.050 4.280 ;
        RECT 273.890 3.670 296.970 4.280 ;
        RECT 297.810 3.670 320.430 4.280 ;
        RECT 321.270 3.670 344.350 4.280 ;
        RECT 345.190 3.670 368.270 4.280 ;
        RECT 369.110 3.670 392.190 4.280 ;
        RECT 393.030 3.670 415.650 4.280 ;
        RECT 416.490 3.670 439.570 4.280 ;
        RECT 440.410 3.670 463.490 4.280 ;
        RECT 464.330 3.670 487.410 4.280 ;
        RECT 488.250 3.670 491.650 4.280 ;
      LAYER met3 ;
        RECT 4.000 489.920 495.600 490.785 ;
        RECT 4.000 483.840 496.000 489.920 ;
        RECT 4.400 482.440 496.000 483.840 ;
        RECT 4.000 474.320 496.000 482.440 ;
        RECT 4.000 472.920 495.600 474.320 ;
        RECT 4.000 456.640 496.000 472.920 ;
        RECT 4.000 455.240 495.600 456.640 ;
        RECT 4.000 450.520 496.000 455.240 ;
        RECT 4.400 449.120 496.000 450.520 ;
        RECT 4.000 439.640 496.000 449.120 ;
        RECT 4.000 438.240 495.600 439.640 ;
        RECT 4.000 422.640 496.000 438.240 ;
        RECT 4.000 421.240 495.600 422.640 ;
        RECT 4.000 417.200 496.000 421.240 ;
        RECT 4.400 415.800 496.000 417.200 ;
        RECT 4.000 404.960 496.000 415.800 ;
        RECT 4.000 403.560 495.600 404.960 ;
        RECT 4.000 387.960 496.000 403.560 ;
        RECT 4.000 386.560 495.600 387.960 ;
        RECT 4.000 383.880 496.000 386.560 ;
        RECT 4.400 382.480 496.000 383.880 ;
        RECT 4.000 370.960 496.000 382.480 ;
        RECT 4.000 369.560 495.600 370.960 ;
        RECT 4.000 353.280 496.000 369.560 ;
        RECT 4.000 351.880 495.600 353.280 ;
        RECT 4.000 350.560 496.000 351.880 ;
        RECT 4.400 349.160 496.000 350.560 ;
        RECT 4.000 336.280 496.000 349.160 ;
        RECT 4.000 334.880 495.600 336.280 ;
        RECT 4.000 319.280 496.000 334.880 ;
        RECT 4.000 317.880 495.600 319.280 ;
        RECT 4.000 317.240 496.000 317.880 ;
        RECT 4.400 315.840 496.000 317.240 ;
        RECT 4.000 301.600 496.000 315.840 ;
        RECT 4.000 300.200 495.600 301.600 ;
        RECT 4.000 284.600 496.000 300.200 ;
        RECT 4.000 283.920 495.600 284.600 ;
        RECT 4.400 283.200 495.600 283.920 ;
        RECT 4.400 282.520 496.000 283.200 ;
        RECT 4.000 267.600 496.000 282.520 ;
        RECT 4.000 266.200 495.600 267.600 ;
        RECT 4.000 250.600 496.000 266.200 ;
        RECT 4.400 249.920 496.000 250.600 ;
        RECT 4.400 249.200 495.600 249.920 ;
        RECT 4.000 248.520 495.600 249.200 ;
        RECT 4.000 232.920 496.000 248.520 ;
        RECT 4.000 231.520 495.600 232.920 ;
        RECT 4.000 217.280 496.000 231.520 ;
        RECT 4.400 215.920 496.000 217.280 ;
        RECT 4.400 215.880 495.600 215.920 ;
        RECT 4.000 214.520 495.600 215.880 ;
        RECT 4.000 198.240 496.000 214.520 ;
        RECT 4.000 196.840 495.600 198.240 ;
        RECT 4.000 183.960 496.000 196.840 ;
        RECT 4.400 182.560 496.000 183.960 ;
        RECT 4.000 181.240 496.000 182.560 ;
        RECT 4.000 179.840 495.600 181.240 ;
        RECT 4.000 164.240 496.000 179.840 ;
        RECT 4.000 162.840 495.600 164.240 ;
        RECT 4.000 150.640 496.000 162.840 ;
        RECT 4.400 149.240 496.000 150.640 ;
        RECT 4.000 146.560 496.000 149.240 ;
        RECT 4.000 145.160 495.600 146.560 ;
        RECT 4.000 129.560 496.000 145.160 ;
        RECT 4.000 128.160 495.600 129.560 ;
        RECT 4.000 117.320 496.000 128.160 ;
        RECT 4.400 115.920 496.000 117.320 ;
        RECT 4.000 112.560 496.000 115.920 ;
        RECT 4.000 111.160 495.600 112.560 ;
        RECT 4.000 94.880 496.000 111.160 ;
        RECT 4.000 93.480 495.600 94.880 ;
        RECT 4.000 84.000 496.000 93.480 ;
        RECT 4.400 82.600 496.000 84.000 ;
        RECT 4.000 77.880 496.000 82.600 ;
        RECT 4.000 76.480 495.600 77.880 ;
        RECT 4.000 60.880 496.000 76.480 ;
        RECT 4.000 59.480 495.600 60.880 ;
        RECT 4.000 50.680 496.000 59.480 ;
        RECT 4.400 49.280 496.000 50.680 ;
        RECT 4.000 43.200 496.000 49.280 ;
        RECT 4.000 41.800 495.600 43.200 ;
        RECT 4.000 26.200 496.000 41.800 ;
        RECT 4.000 24.800 495.600 26.200 ;
        RECT 4.000 17.360 496.000 24.800 ;
        RECT 4.400 15.960 496.000 17.360 ;
        RECT 4.000 9.200 496.000 15.960 ;
        RECT 4.000 8.335 495.600 9.200 ;
      LAYER met4 ;
        RECT 230.295 13.095 251.040 485.345 ;
        RECT 253.440 13.095 327.840 485.345 ;
        RECT 330.240 13.095 404.640 485.345 ;
        RECT 407.040 13.095 454.185 485.345 ;
  END
END Motor_Top
END LIBRARY

