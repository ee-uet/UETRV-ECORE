magic
tech sky130A
magscale 1 2
timestamp 1647892870
<< metal1 >>
rect 204254 325660 204260 325712
rect 204312 325700 204318 325712
rect 207014 325700 207020 325712
rect 204312 325672 207020 325700
rect 204312 325660 204318 325672
rect 207014 325660 207020 325672
rect 207072 325660 207078 325712
rect 193214 306348 193220 306400
rect 193272 306388 193278 306400
rect 207014 306388 207020 306400
rect 193272 306360 207020 306388
rect 193272 306348 193278 306360
rect 207014 306348 207020 306360
rect 207072 306348 207078 306400
rect 190454 304988 190460 305040
rect 190512 305028 190518 305040
rect 207014 305028 207020 305040
rect 190512 305000 207020 305028
rect 190512 304988 190518 305000
rect 207014 304988 207020 305000
rect 207072 304988 207078 305040
rect 67818 298256 67824 298308
rect 67876 298296 67882 298308
rect 227714 298296 227720 298308
rect 67876 298268 227720 298296
rect 67876 298256 67882 298268
rect 227714 298256 227720 298268
rect 227772 298256 227778 298308
rect 69290 298188 69296 298240
rect 69348 298228 69354 298240
rect 229094 298228 229100 298240
rect 69348 298200 229100 298228
rect 69348 298188 69354 298200
rect 229094 298188 229100 298200
rect 229152 298188 229158 298240
rect 55214 298120 55220 298172
rect 55272 298160 55278 298172
rect 55858 298160 55864 298172
rect 55272 298132 55864 298160
rect 55272 298120 55278 298132
rect 55858 298120 55864 298132
rect 55916 298160 55922 298172
rect 215846 298160 215852 298172
rect 55916 298132 215852 298160
rect 55916 298120 55922 298132
rect 215846 298120 215852 298132
rect 215904 298120 215910 298172
rect 76834 297984 76840 298036
rect 76892 298024 76898 298036
rect 79318 298024 79324 298036
rect 76892 297996 79324 298024
rect 76892 297984 76898 297996
rect 79318 297984 79324 297996
rect 79376 297984 79382 298036
rect 97074 297440 97080 297492
rect 97132 297480 97138 297492
rect 130470 297480 130476 297492
rect 97132 297452 130476 297480
rect 97132 297440 97138 297452
rect 130470 297440 130476 297452
rect 130528 297440 130534 297492
rect 89162 297372 89168 297424
rect 89220 297412 89226 297424
rect 130378 297412 130384 297424
rect 89220 297384 130384 297412
rect 89220 297372 89226 297384
rect 130378 297372 130384 297384
rect 130436 297372 130442 297424
rect 75546 297304 75552 297356
rect 75604 297344 75610 297356
rect 131758 297344 131764 297356
rect 75604 297316 131764 297344
rect 75604 297304 75610 297316
rect 131758 297304 131764 297316
rect 131816 297304 131822 297356
rect 70210 297236 70216 297288
rect 70268 297276 70274 297288
rect 229278 297276 229284 297288
rect 70268 297248 229284 297276
rect 70268 297236 70274 297248
rect 229278 297236 229284 297248
rect 229336 297236 229342 297288
rect 106642 297168 106648 297220
rect 106700 297208 106706 297220
rect 341518 297208 341524 297220
rect 106700 297180 341524 297208
rect 106700 297168 106706 297180
rect 341518 297168 341524 297180
rect 341576 297168 341582 297220
rect 107746 297100 107752 297152
rect 107804 297140 107810 297152
rect 345658 297140 345664 297152
rect 107804 297112 345664 297140
rect 107804 297100 107810 297112
rect 345658 297100 345664 297112
rect 345716 297100 345722 297152
rect 111610 297032 111616 297084
rect 111668 297072 111674 297084
rect 409046 297072 409052 297084
rect 111668 297044 409052 297072
rect 111668 297032 111674 297044
rect 409046 297032 409052 297044
rect 409104 297032 409110 297084
rect 105538 296964 105544 297016
rect 105596 297004 105602 297016
rect 408862 297004 408868 297016
rect 105596 296976 408868 297004
rect 105596 296964 105602 296976
rect 408862 296964 408868 296976
rect 408920 296964 408926 297016
rect 104250 296896 104256 296948
rect 104308 296936 104314 296948
rect 409322 296936 409328 296948
rect 104308 296908 409328 296936
rect 104308 296896 104314 296908
rect 409322 296896 409328 296908
rect 409380 296896 409386 296948
rect 102962 296828 102968 296880
rect 103020 296868 103026 296880
rect 409230 296868 409236 296880
rect 103020 296840 409236 296868
rect 103020 296828 103026 296840
rect 409230 296828 409236 296840
rect 409288 296828 409294 296880
rect 102042 296760 102048 296812
rect 102100 296800 102106 296812
rect 409138 296800 409144 296812
rect 102100 296772 409144 296800
rect 102100 296760 102106 296772
rect 409138 296760 409144 296772
rect 409196 296760 409202 296812
rect 65794 296692 65800 296744
rect 65852 296732 65858 296744
rect 408954 296732 408960 296744
rect 65852 296704 408960 296732
rect 65852 296692 65858 296704
rect 408954 296692 408960 296704
rect 409012 296692 409018 296744
rect 234614 295944 234620 295996
rect 234672 295984 234678 295996
rect 242894 295984 242900 295996
rect 234672 295956 242900 295984
rect 234672 295944 234678 295956
rect 242894 295944 242900 295956
rect 242952 295944 242958 295996
rect 49418 291796 49424 291848
rect 49476 291836 49482 291848
rect 371234 291836 371240 291848
rect 49476 291808 371240 291836
rect 49476 291796 49482 291808
rect 371234 291796 371240 291808
rect 371292 291796 371298 291848
rect 47762 287648 47768 287700
rect 47820 287688 47826 287700
rect 409966 287688 409972 287700
rect 47820 287660 409972 287688
rect 47820 287648 47826 287660
rect 409966 287648 409972 287660
rect 410024 287648 410030 287700
rect 208118 282344 208124 282396
rect 208176 282384 208182 282396
rect 213914 282384 213920 282396
rect 208176 282356 213920 282384
rect 208176 282344 208182 282356
rect 213914 282344 213920 282356
rect 213972 282344 213978 282396
rect 194594 282276 194600 282328
rect 194652 282316 194658 282328
rect 224954 282316 224960 282328
rect 194652 282288 224960 282316
rect 194652 282276 194658 282288
rect 224954 282276 224960 282288
rect 225012 282276 225018 282328
rect 266170 282276 266176 282328
rect 266228 282316 266234 282328
rect 358814 282316 358820 282328
rect 266228 282288 358820 282316
rect 266228 282276 266234 282288
rect 358814 282276 358820 282288
rect 358872 282276 358878 282328
rect 197354 282208 197360 282260
rect 197412 282248 197418 282260
rect 237374 282248 237380 282260
rect 197412 282220 237380 282248
rect 197412 282208 197418 282220
rect 237374 282208 237380 282220
rect 237432 282208 237438 282260
rect 267458 282208 267464 282260
rect 267516 282248 267522 282260
rect 364334 282248 364340 282260
rect 267516 282220 364340 282248
rect 267516 282208 267522 282220
rect 364334 282208 364340 282220
rect 364392 282208 364398 282260
rect 47854 282140 47860 282192
rect 47912 282180 47918 282192
rect 410058 282180 410064 282192
rect 47912 282152 410064 282180
rect 47912 282140 47918 282152
rect 410058 282140 410064 282152
rect 410116 282140 410122 282192
rect 218054 280848 218060 280900
rect 218112 280888 218118 280900
rect 229094 280888 229100 280900
rect 218112 280860 229100 280888
rect 218112 280848 218118 280860
rect 229094 280848 229100 280860
rect 229152 280848 229158 280900
rect 209590 280780 209596 280832
rect 209648 280820 209654 280832
rect 231854 280820 231860 280832
rect 209648 280792 231860 280820
rect 209648 280780 209654 280792
rect 231854 280780 231860 280792
rect 231912 280780 231918 280832
rect 248230 280780 248236 280832
rect 248288 280820 248294 280832
rect 259454 280820 259460 280832
rect 248288 280792 259460 280820
rect 248288 280780 248294 280792
rect 259454 280780 259460 280792
rect 259512 280780 259518 280832
rect 209498 279624 209504 279676
rect 209556 279664 209562 279676
rect 222194 279664 222200 279676
rect 209556 279636 222200 279664
rect 209556 279624 209562 279636
rect 222194 279624 222200 279636
rect 222252 279624 222258 279676
rect 85298 279556 85304 279608
rect 85356 279596 85362 279608
rect 389174 279596 389180 279608
rect 85356 279568 389180 279596
rect 85356 279556 85362 279568
rect 389174 279556 389180 279568
rect 389232 279556 389238 279608
rect 49510 279488 49516 279540
rect 49568 279528 49574 279540
rect 373994 279528 374000 279540
rect 49568 279500 374000 279528
rect 49568 279488 49574 279500
rect 373994 279488 374000 279500
rect 374052 279488 374058 279540
rect 47670 279420 47676 279472
rect 47728 279460 47734 279472
rect 409874 279460 409880 279472
rect 47728 279432 409880 279460
rect 47728 279420 47734 279432
rect 409874 279420 409880 279432
rect 409932 279420 409938 279472
rect 245562 273912 245568 273964
rect 245620 273952 245626 273964
rect 280154 273952 280160 273964
rect 245620 273924 280160 273952
rect 245620 273912 245626 273924
rect 280154 273912 280160 273924
rect 280212 273912 280218 273964
rect 246758 271804 246764 271856
rect 246816 271844 246822 271856
rect 248414 271844 248420 271856
rect 246816 271816 248420 271844
rect 246816 271804 246822 271816
rect 248414 271804 248420 271816
rect 248472 271804 248478 271856
rect 264790 268404 264796 268456
rect 264848 268444 264854 268456
rect 354674 268444 354680 268456
rect 264848 268416 354680 268444
rect 264848 268404 264854 268416
rect 354674 268404 354680 268416
rect 354732 268404 354738 268456
rect 242802 268336 242808 268388
rect 242860 268376 242866 268388
rect 266354 268376 266360 268388
rect 242860 268348 266360 268376
rect 242860 268336 242866 268348
rect 266354 268336 266360 268348
rect 266412 268336 266418 268388
rect 267550 268336 267556 268388
rect 267608 268376 267614 268388
rect 368474 268376 368480 268388
rect 267608 268348 368480 268376
rect 267608 268336 267614 268348
rect 368474 268336 368480 268348
rect 368532 268336 368538 268388
rect 229094 268132 229100 268184
rect 229152 268172 229158 268184
rect 234706 268172 234712 268184
rect 229152 268144 234712 268172
rect 229152 268132 229158 268144
rect 234706 268132 234712 268144
rect 234764 268132 234770 268184
rect 260650 267112 260656 267164
rect 260708 267152 260714 267164
rect 341058 267152 341064 267164
rect 260708 267124 341064 267152
rect 260708 267112 260714 267124
rect 341058 267112 341064 267124
rect 341116 267112 341122 267164
rect 262030 267044 262036 267096
rect 262088 267084 262094 267096
rect 345566 267084 345572 267096
rect 262088 267056 345572 267084
rect 262088 267044 262094 267056
rect 345566 267044 345572 267056
rect 345624 267044 345630 267096
rect 263410 266976 263416 267028
rect 263468 267016 263474 267028
rect 350534 267016 350540 267028
rect 263468 266988 350540 267016
rect 263468 266976 263474 266988
rect 350534 266976 350540 266988
rect 350592 266976 350598 267028
rect 257798 265752 257804 265804
rect 257856 265792 257862 265804
rect 327258 265792 327264 265804
rect 257856 265764 327264 265792
rect 257856 265752 257862 265764
rect 327258 265752 327264 265764
rect 327316 265752 327322 265804
rect 259270 265684 259276 265736
rect 259328 265724 259334 265736
rect 331858 265724 331864 265736
rect 259328 265696 331864 265724
rect 259328 265684 259334 265696
rect 331858 265684 331864 265696
rect 331916 265684 331922 265736
rect 259178 265616 259184 265668
rect 259236 265656 259242 265668
rect 336734 265656 336740 265668
rect 259236 265628 336740 265656
rect 259236 265616 259242 265628
rect 336734 265616 336740 265628
rect 336792 265616 336798 265668
rect 253750 264392 253756 264444
rect 253808 264432 253814 264444
rect 313274 264432 313280 264444
rect 253808 264404 313280 264432
rect 253808 264392 253814 264404
rect 313274 264392 313280 264404
rect 313332 264392 313338 264444
rect 255130 264324 255136 264376
rect 255188 264364 255194 264376
rect 318058 264364 318064 264376
rect 255188 264336 318064 264364
rect 255188 264324 255194 264336
rect 318058 264324 318064 264336
rect 318116 264324 318122 264376
rect 256510 264256 256516 264308
rect 256568 264296 256574 264308
rect 322934 264296 322940 264308
rect 256568 264268 322940 264296
rect 256568 264256 256574 264268
rect 322934 264256 322940 264268
rect 322992 264256 322998 264308
rect 100570 264188 100576 264240
rect 100628 264228 100634 264240
rect 399018 264228 399024 264240
rect 100628 264200 399024 264228
rect 100628 264188 100634 264200
rect 399018 264188 399024 264200
rect 399076 264188 399082 264240
rect 248322 263100 248328 263152
rect 248380 263140 248386 263152
rect 290274 263140 290280 263152
rect 248380 263112 290280 263140
rect 248380 263100 248386 263112
rect 290274 263100 290280 263112
rect 290332 263100 290338 263152
rect 252278 263032 252284 263084
rect 252336 263072 252342 263084
rect 304074 263072 304080 263084
rect 252336 263044 304080 263072
rect 252336 263032 252342 263044
rect 304074 263032 304080 263044
rect 304132 263032 304138 263084
rect 252370 262964 252376 263016
rect 252428 263004 252434 263016
rect 309226 263004 309232 263016
rect 252428 262976 309232 263004
rect 252428 262964 252434 262976
rect 309226 262964 309232 262976
rect 309284 262964 309290 263016
rect 96430 262896 96436 262948
rect 96488 262936 96494 262948
rect 411898 262936 411904 262948
rect 96488 262908 411904 262936
rect 96488 262896 96494 262908
rect 411898 262896 411904 262908
rect 411956 262896 411962 262948
rect 81250 262828 81256 262880
rect 81308 262868 81314 262880
rect 411530 262868 411536 262880
rect 81308 262840 411536 262868
rect 81308 262828 81314 262840
rect 411530 262828 411536 262840
rect 411588 262828 411594 262880
rect 255222 261808 255228 261860
rect 255280 261848 255286 261860
rect 283282 261848 283288 261860
rect 255280 261820 283288 261848
rect 255280 261808 255286 261820
rect 283282 261808 283288 261820
rect 283340 261808 283346 261860
rect 256602 261740 256608 261792
rect 256660 261780 256666 261792
rect 287882 261780 287888 261792
rect 256660 261752 287888 261780
rect 256660 261740 256666 261752
rect 287882 261740 287888 261752
rect 287940 261740 287946 261792
rect 211522 261672 211528 261724
rect 211580 261712 211586 261724
rect 231946 261712 231952 261724
rect 211580 261684 231952 261712
rect 211580 261672 211586 261684
rect 231946 261672 231952 261684
rect 232004 261672 232010 261724
rect 246850 261672 246856 261724
rect 246908 261712 246914 261724
rect 255498 261712 255504 261724
rect 246908 261684 255504 261712
rect 246908 261672 246914 261684
rect 255498 261672 255504 261684
rect 255556 261672 255562 261724
rect 259362 261672 259368 261724
rect 259420 261712 259426 261724
rect 302326 261712 302332 261724
rect 259420 261684 302332 261712
rect 259420 261672 259426 261684
rect 302326 261672 302332 261684
rect 302384 261672 302390 261724
rect 88150 261604 88156 261656
rect 88208 261644 88214 261656
rect 387794 261644 387800 261656
rect 88208 261616 387800 261644
rect 88208 261604 88214 261616
rect 387794 261604 387800 261616
rect 387852 261604 387858 261656
rect 90910 261536 90916 261588
rect 90968 261576 90974 261588
rect 392026 261576 392032 261588
rect 90968 261548 392032 261576
rect 90968 261536 90974 261548
rect 392026 261536 392032 261548
rect 392084 261536 392090 261588
rect 86678 261468 86684 261520
rect 86736 261508 86742 261520
rect 411622 261508 411628 261520
rect 86736 261480 411628 261508
rect 86736 261468 86742 261480
rect 411622 261468 411628 261480
rect 411680 261468 411686 261520
rect 252462 260448 252468 260500
rect 252520 260488 252526 260500
rect 274082 260488 274088 260500
rect 252520 260460 274088 260488
rect 252520 260448 252526 260460
rect 274082 260448 274088 260460
rect 274140 260448 274146 260500
rect 225322 260380 225328 260432
rect 225380 260420 225386 260432
rect 241514 260420 241520 260432
rect 225380 260392 241520 260420
rect 225380 260380 225386 260392
rect 241514 260380 241520 260392
rect 241572 260380 241578 260432
rect 253842 260380 253848 260432
rect 253900 260420 253906 260432
rect 278774 260420 278780 260432
rect 253900 260392 278780 260420
rect 253900 260380 253906 260392
rect 278774 260380 278780 260392
rect 278832 260380 278838 260432
rect 74442 260312 74448 260364
rect 74500 260352 74506 260364
rect 148318 260352 148324 260364
rect 74500 260324 148324 260352
rect 74500 260312 74506 260324
rect 148318 260312 148324 260324
rect 148376 260312 148382 260364
rect 216122 260312 216128 260364
rect 216180 260352 216186 260364
rect 240134 260352 240140 260364
rect 216180 260324 240140 260352
rect 216180 260312 216186 260324
rect 240134 260312 240140 260324
rect 240192 260312 240198 260364
rect 273070 260312 273076 260364
rect 273128 260352 273134 260364
rect 348050 260352 348056 260364
rect 273128 260324 348056 260352
rect 273128 260312 273134 260324
rect 348050 260312 348056 260324
rect 348108 260312 348114 260364
rect 79870 260244 79876 260296
rect 79928 260284 79934 260296
rect 153194 260284 153200 260296
rect 79928 260256 153200 260284
rect 79928 260244 79934 260256
rect 153194 260244 153200 260256
rect 153252 260244 153258 260296
rect 202138 260244 202144 260296
rect 202196 260284 202202 260296
rect 230474 260284 230480 260296
rect 202196 260256 230480 260284
rect 202196 260244 202202 260256
rect 230474 260244 230480 260256
rect 230532 260244 230538 260296
rect 237190 260244 237196 260296
rect 237248 260284 237254 260296
rect 244366 260284 244372 260296
rect 237248 260256 244372 260284
rect 237248 260244 237254 260256
rect 244366 260244 244372 260256
rect 244424 260244 244430 260296
rect 250990 260244 250996 260296
rect 251048 260284 251054 260296
rect 269298 260284 269304 260296
rect 251048 260256 269304 260284
rect 251048 260244 251054 260256
rect 269298 260244 269304 260256
rect 269356 260244 269362 260296
rect 273162 260244 273168 260296
rect 273220 260284 273226 260296
rect 352650 260284 352656 260296
rect 273220 260256 352656 260284
rect 273220 260244 273226 260256
rect 352650 260244 352656 260256
rect 352708 260244 352714 260296
rect 115842 260176 115848 260228
rect 115900 260216 115906 260228
rect 403618 260216 403624 260228
rect 115900 260188 403624 260216
rect 115900 260176 115906 260188
rect 403618 260176 403624 260188
rect 403676 260176 403682 260228
rect 112990 260108 112996 260160
rect 113048 260148 113054 260160
rect 401594 260148 401600 260160
rect 113048 260120 401600 260148
rect 113048 260108 113054 260120
rect 401594 260108 401600 260120
rect 401652 260108 401658 260160
rect 241606 260040 241612 260092
rect 241664 260080 241670 260092
rect 244274 260080 244280 260092
rect 241664 260052 244280 260080
rect 241664 260040 241670 260052
rect 244274 260040 244280 260052
rect 244332 260040 244338 260092
rect 244090 258952 244096 259004
rect 244148 258992 244154 259004
rect 276290 258992 276296 259004
rect 244148 258964 276296 258992
rect 244148 258952 244154 258964
rect 276290 258952 276296 258964
rect 276348 258952 276354 259004
rect 249610 258884 249616 258936
rect 249668 258924 249674 258936
rect 294874 258924 294880 258936
rect 249668 258896 294880 258924
rect 249668 258884 249674 258896
rect 294874 258884 294880 258896
rect 294932 258884 294938 258936
rect 251082 258816 251088 258868
rect 251140 258856 251146 258868
rect 299474 258856 299480 258868
rect 251140 258828 299480 258856
rect 251140 258816 251146 258828
rect 299474 258816 299480 258828
rect 299532 258816 299538 258868
rect 93578 258748 93584 258800
rect 93636 258788 93642 258800
rect 410242 258788 410248 258800
rect 93636 258760 410248 258788
rect 93636 258748 93642 258760
rect 410242 258748 410248 258760
rect 410300 258748 410306 258800
rect 85390 258680 85396 258732
rect 85448 258720 85454 258732
rect 411346 258720 411352 258732
rect 85448 258692 411352 258720
rect 85448 258680 85454 258692
rect 411346 258680 411352 258692
rect 411404 258680 411410 258732
rect 246942 257660 246948 257712
rect 247000 257700 247006 257712
rect 285674 257700 285680 257712
rect 247000 257672 285680 257700
rect 247000 257660 247006 257672
rect 285674 257660 285680 257672
rect 285732 257660 285738 257712
rect 260742 257592 260748 257644
rect 260800 257632 260806 257644
rect 306558 257632 306564 257644
rect 260800 257604 306564 257632
rect 260800 257592 260806 257604
rect 306558 257592 306564 257604
rect 306616 257592 306622 257644
rect 244182 257524 244188 257576
rect 244240 257564 244246 257576
rect 271874 257564 271880 257576
rect 244240 257536 271880 257564
rect 244240 257524 244246 257536
rect 271874 257524 271880 257536
rect 271932 257524 271938 257576
rect 277302 257524 277308 257576
rect 277360 257564 277366 257576
rect 366726 257564 366732 257576
rect 277360 257536 366732 257564
rect 277360 257524 277366 257536
rect 366726 257524 366732 257536
rect 366784 257524 366790 257576
rect 108850 257456 108856 257508
rect 108908 257496 108914 257508
rect 396718 257496 396724 257508
rect 108908 257468 396724 257496
rect 108908 257456 108914 257468
rect 396718 257456 396724 257468
rect 396776 257456 396782 257508
rect 104710 257388 104716 257440
rect 104768 257428 104774 257440
rect 394694 257428 394700 257440
rect 104768 257400 394700 257428
rect 104768 257388 104774 257400
rect 394694 257388 394700 257400
rect 394752 257388 394758 257440
rect 81342 257320 81348 257372
rect 81400 257360 81406 257372
rect 375926 257360 375932 257372
rect 81400 257332 375932 257360
rect 81400 257320 81406 257332
rect 375926 257320 375932 257332
rect 375984 257320 375990 257372
rect 221458 256232 221464 256284
rect 221516 256272 221522 256284
rect 233234 256272 233240 256284
rect 221516 256244 233240 256272
rect 221516 256232 221522 256244
rect 233234 256232 233240 256244
rect 233292 256232 233298 256284
rect 257890 256232 257896 256284
rect 257948 256272 257954 256284
rect 297174 256272 297180 256284
rect 257948 256244 297180 256272
rect 257948 256232 257954 256244
rect 297174 256232 297180 256244
rect 297232 256232 297238 256284
rect 209498 256164 209504 256216
rect 209556 256204 209562 256216
rect 227714 256204 227720 256216
rect 209556 256176 227720 256204
rect 209556 256164 209562 256176
rect 227714 256164 227720 256176
rect 227772 256164 227778 256216
rect 262122 256164 262128 256216
rect 262180 256204 262186 256216
rect 311158 256204 311164 256216
rect 262180 256176 311164 256204
rect 262180 256164 262186 256176
rect 311158 256164 311164 256176
rect 311216 256164 311222 256216
rect 201402 256096 201408 256148
rect 201460 256136 201466 256148
rect 226334 256136 226340 256148
rect 201460 256108 226340 256136
rect 201460 256096 201466 256108
rect 226334 256096 226340 256108
rect 226392 256096 226398 256148
rect 263502 256096 263508 256148
rect 263560 256136 263566 256148
rect 316034 256136 316040 256148
rect 263560 256108 316040 256136
rect 263560 256096 263566 256108
rect 316034 256096 316040 256108
rect 316092 256096 316098 256148
rect 97810 256028 97816 256080
rect 97868 256068 97874 256080
rect 410426 256068 410432 256080
rect 97868 256040 410432 256068
rect 97868 256028 97874 256040
rect 410426 256028 410432 256040
rect 410484 256028 410490 256080
rect 84010 255960 84016 256012
rect 84068 256000 84074 256012
rect 411438 256000 411444 256012
rect 84068 255972 411444 256000
rect 84068 255960 84074 255972
rect 411438 255960 411444 255972
rect 411496 255960 411502 256012
rect 209682 254736 209688 254788
rect 209740 254776 209746 254788
rect 253198 254776 253204 254788
rect 209740 254748 253204 254776
rect 209740 254736 209746 254748
rect 253198 254736 253204 254748
rect 253256 254736 253262 254788
rect 257982 254736 257988 254788
rect 258040 254776 258046 254788
rect 292574 254776 292580 254788
rect 258040 254748 292580 254776
rect 258040 254736 258046 254748
rect 292574 254736 292580 254748
rect 292632 254736 292638 254788
rect 92290 254668 92296 254720
rect 92348 254708 92354 254720
rect 410334 254708 410340 254720
rect 92348 254680 410340 254708
rect 92348 254668 92354 254680
rect 410334 254668 410340 254680
rect 410392 254668 410398 254720
rect 91002 254600 91008 254652
rect 91060 254640 91066 254652
rect 410150 254640 410156 254652
rect 91060 254612 410156 254640
rect 91060 254600 91066 254612
rect 410150 254600 410156 254612
rect 410208 254600 410214 254652
rect 82630 254532 82636 254584
rect 82688 254572 82694 254584
rect 411254 254572 411260 254584
rect 82688 254544 411260 254572
rect 82688 254532 82694 254544
rect 411254 254532 411260 254544
rect 411312 254532 411318 254584
rect 228450 253852 228456 253904
rect 228508 253892 228514 253904
rect 229186 253892 229192 253904
rect 228508 253864 229192 253892
rect 228508 253852 228514 253864
rect 229186 253852 229192 253864
rect 229244 253852 229250 253904
rect 264882 253648 264888 253700
rect 264940 253688 264946 253700
rect 320358 253688 320364 253700
rect 264940 253660 320364 253688
rect 264940 253648 264946 253660
rect 320358 253648 320364 253660
rect 320416 253648 320422 253700
rect 266262 253580 266268 253632
rect 266320 253620 266326 253632
rect 324958 253620 324964 253632
rect 266320 253592 324964 253620
rect 266320 253580 266326 253592
rect 324958 253580 324964 253592
rect 325016 253580 325022 253632
rect 267642 253512 267648 253564
rect 267700 253552 267706 253564
rect 329834 253552 329840 253564
rect 267700 253524 329840 253552
rect 267700 253512 267706 253524
rect 329834 253512 329840 253524
rect 329892 253512 329898 253564
rect 269022 253444 269028 253496
rect 269080 253484 269086 253496
rect 334342 253484 334348 253496
rect 269080 253456 334348 253484
rect 269080 253444 269086 253456
rect 334342 253444 334348 253456
rect 334400 253444 334406 253496
rect 208210 253376 208216 253428
rect 208268 253416 208274 253428
rect 239398 253416 239404 253428
rect 208268 253388 239404 253416
rect 208268 253376 208274 253388
rect 239398 253376 239404 253388
rect 239456 253376 239462 253428
rect 270402 253376 270408 253428
rect 270460 253416 270466 253428
rect 338942 253416 338948 253428
rect 270460 253388 338948 253416
rect 270460 253376 270466 253388
rect 338942 253376 338948 253388
rect 339000 253376 339006 253428
rect 271782 253308 271788 253360
rect 271840 253348 271846 253360
rect 343634 253348 343640 253360
rect 271840 253320 343640 253348
rect 271840 253308 271846 253320
rect 343634 253308 343640 253320
rect 343692 253308 343698 253360
rect 207658 253240 207664 253292
rect 207716 253280 207722 253292
rect 238754 253280 238760 253292
rect 207716 253252 238760 253280
rect 207716 253240 207722 253252
rect 238754 253240 238760 253252
rect 238812 253240 238818 253292
rect 240042 253240 240048 253292
rect 240100 253280 240106 253292
rect 258074 253280 258080 253292
rect 240100 253252 258080 253280
rect 240100 253240 240106 253252
rect 258074 253240 258080 253252
rect 258132 253240 258138 253292
rect 274542 253240 274548 253292
rect 274600 253280 274606 253292
rect 357526 253280 357532 253292
rect 274600 253252 357532 253280
rect 274600 253240 274606 253252
rect 357526 253240 357532 253252
rect 357584 253240 357590 253292
rect 208302 253172 208308 253224
rect 208360 253212 208366 253224
rect 246390 253212 246396 253224
rect 208360 253184 246396 253212
rect 208360 253172 208366 253184
rect 246390 253172 246396 253184
rect 246448 253172 246454 253224
rect 249702 253172 249708 253224
rect 249760 253212 249766 253224
rect 264974 253212 264980 253224
rect 249760 253184 264980 253212
rect 249760 253172 249766 253184
rect 264974 253172 264980 253184
rect 265032 253172 265038 253224
rect 275922 253172 275928 253224
rect 275980 253212 275986 253224
rect 362126 253212 362132 253224
rect 275980 253184 362132 253212
rect 275980 253172 275986 253184
rect 362126 253172 362132 253184
rect 362184 253172 362190 253224
rect 67542 252492 67548 252544
rect 67600 252532 67606 252544
rect 200390 252532 200396 252544
rect 67600 252504 200396 252532
rect 67600 252492 67606 252504
rect 200390 252492 200396 252504
rect 200448 252532 200454 252544
rect 201402 252532 201408 252544
rect 200448 252504 201408 252532
rect 200448 252492 200454 252504
rect 201402 252492 201408 252504
rect 201460 252492 201466 252544
rect 238662 252152 238668 252204
rect 238720 252192 238726 252204
rect 251174 252192 251180 252204
rect 238720 252164 251180 252192
rect 238720 252152 238726 252164
rect 251174 252152 251180 252164
rect 251232 252152 251238 252204
rect 345658 252152 345664 252204
rect 345716 252192 345722 252204
rect 408494 252192 408500 252204
rect 345716 252164 408500 252192
rect 345716 252152 345722 252164
rect 408494 252152 408500 252164
rect 408552 252152 408558 252204
rect 241422 252084 241428 252136
rect 241480 252124 241486 252136
rect 262582 252124 262588 252136
rect 241480 252096 262588 252124
rect 241480 252084 241486 252096
rect 262582 252084 262588 252096
rect 262640 252084 262646 252136
rect 341518 252084 341524 252136
rect 341576 252124 341582 252136
rect 406102 252124 406108 252136
rect 341576 252096 406108 252124
rect 341576 252084 341582 252096
rect 406102 252084 406108 252096
rect 406160 252084 406166 252136
rect 148318 252016 148324 252068
rect 148376 252056 148382 252068
rect 378318 252056 378324 252068
rect 148376 252028 378324 252056
rect 148376 252016 148382 252028
rect 378318 252016 378324 252028
rect 378376 252016 378382 252068
rect 153194 251948 153200 252000
rect 153252 251988 153258 252000
rect 385310 251988 385316 252000
rect 153252 251960 385316 251988
rect 153252 251948 153258 251960
rect 385310 251948 385316 251960
rect 385368 251948 385374 252000
rect 79318 251880 79324 251932
rect 79376 251920 79382 251932
rect 380986 251920 380992 251932
rect 79376 251892 380992 251920
rect 79376 251880 79382 251892
rect 380986 251880 380992 251892
rect 381044 251880 381050 251932
rect 77110 251812 77116 251864
rect 77168 251852 77174 251864
rect 382918 251852 382924 251864
rect 77168 251824 382924 251852
rect 77168 251812 77174 251824
rect 382918 251812 382924 251824
rect 382976 251812 382982 251864
rect 101950 250588 101956 250640
rect 102008 250628 102014 250640
rect 410518 250628 410524 250640
rect 102008 250600 410524 250628
rect 102008 250588 102014 250600
rect 410518 250588 410524 250600
rect 410576 250588 410582 250640
rect 82722 250520 82728 250572
rect 82780 250560 82786 250572
rect 411806 250560 411812 250572
rect 82780 250532 411812 250560
rect 82780 250520 82786 250532
rect 411806 250520 411812 250532
rect 411864 250520 411870 250572
rect 78490 250452 78496 250504
rect 78548 250492 78554 250504
rect 411714 250492 411720 250504
rect 78548 250464 411720 250492
rect 78548 250452 78554 250464
rect 411714 250452 411720 250464
rect 411772 250452 411778 250504
rect 114462 249704 114468 249756
rect 114520 249744 114526 249756
rect 186314 249744 186320 249756
rect 114520 249716 186320 249744
rect 114520 249704 114526 249716
rect 186314 249704 186320 249716
rect 186372 249704 186378 249756
rect 106090 248344 106096 248396
rect 106148 248384 106154 248396
rect 186406 248384 186412 248396
rect 106148 248356 186412 248384
rect 106148 248344 106154 248356
rect 186406 248344 186412 248356
rect 186464 248344 186470 248396
rect 107470 248276 107476 248328
rect 107528 248316 107534 248328
rect 186314 248316 186320 248328
rect 107528 248288 186320 248316
rect 107528 248276 107534 248288
rect 186314 248276 186320 248288
rect 186372 248276 186378 248328
rect 95050 246984 95056 247036
rect 95108 247024 95114 247036
rect 186314 247024 186320 247036
rect 95108 246996 186320 247024
rect 95108 246984 95114 246996
rect 186314 246984 186320 246996
rect 186372 246984 186378 247036
rect 85482 246304 85488 246356
rect 85540 246344 85546 246356
rect 187142 246344 187148 246356
rect 85540 246316 187148 246344
rect 85540 246304 85546 246316
rect 187142 246304 187148 246316
rect 187200 246304 187206 246356
rect 103330 245556 103336 245608
rect 103388 245596 103394 245608
rect 186314 245596 186320 245608
rect 103388 245568 186320 245596
rect 103388 245556 103394 245568
rect 186314 245556 186320 245568
rect 186372 245556 186378 245608
rect 101858 244196 101864 244248
rect 101916 244236 101922 244248
rect 186314 244236 186320 244248
rect 101916 244208 186320 244236
rect 101916 244196 101922 244208
rect 186314 244196 186320 244208
rect 186372 244196 186378 244248
rect 100662 242836 100668 242888
rect 100720 242876 100726 242888
rect 186314 242876 186320 242888
rect 100720 242848 186320 242876
rect 100720 242836 100726 242848
rect 186314 242836 186320 242848
rect 186372 242836 186378 242888
rect 88242 241408 88248 241460
rect 88300 241448 88306 241460
rect 186314 241448 186320 241460
rect 88300 241420 186320 241448
rect 88300 241408 88306 241420
rect 186314 241408 186320 241420
rect 186372 241408 186378 241460
rect 95142 240048 95148 240100
rect 95200 240088 95206 240100
rect 186406 240088 186412 240100
rect 95200 240060 186412 240088
rect 95200 240048 95206 240060
rect 186406 240048 186412 240060
rect 186464 240048 186470 240100
rect 96522 239980 96528 240032
rect 96580 240020 96586 240032
rect 186314 240020 186320 240032
rect 96580 239992 186320 240020
rect 96580 239980 96586 239992
rect 186314 239980 186320 239992
rect 186372 239980 186378 240032
rect 84102 237328 84108 237380
rect 84160 237368 84166 237380
rect 186314 237368 186320 237380
rect 84160 237340 186320 237368
rect 84160 237328 84166 237340
rect 186314 237328 186320 237340
rect 186372 237328 186378 237380
rect 89530 235900 89536 235952
rect 89588 235940 89594 235952
rect 186314 235940 186320 235952
rect 89588 235912 186320 235940
rect 89588 235900 89594 235912
rect 186314 235900 186320 235912
rect 186372 235900 186378 235952
rect 86770 234540 86776 234592
rect 86828 234580 86834 234592
rect 186314 234580 186320 234592
rect 86828 234552 186320 234580
rect 86828 234540 86834 234552
rect 186314 234540 186320 234552
rect 186372 234540 186378 234592
rect 49602 233180 49608 233232
rect 49660 233220 49666 233232
rect 186406 233220 186412 233232
rect 49660 233192 186412 233220
rect 49660 233180 49666 233192
rect 186406 233180 186412 233192
rect 186464 233180 186470 233232
rect 86862 233112 86868 233164
rect 86920 233152 86926 233164
rect 186314 233152 186320 233164
rect 86920 233124 186320 233152
rect 86920 233112 86926 233124
rect 186314 233112 186320 233124
rect 186372 233112 186378 233164
rect 73062 231752 73068 231804
rect 73120 231792 73126 231804
rect 186314 231792 186320 231804
rect 73120 231764 186320 231792
rect 73120 231752 73126 231764
rect 186314 231752 186320 231764
rect 186372 231752 186378 231804
rect 71682 230392 71688 230444
rect 71740 230432 71746 230444
rect 186314 230432 186320 230444
rect 71740 230404 186320 230432
rect 71740 230392 71746 230404
rect 186314 230392 186320 230404
rect 186372 230392 186378 230444
rect 169018 227740 169024 227792
rect 169076 227780 169082 227792
rect 186314 227780 186320 227792
rect 169076 227752 186320 227780
rect 169076 227740 169082 227752
rect 186314 227740 186320 227752
rect 186372 227740 186378 227792
rect 148318 226312 148324 226364
rect 148376 226352 148382 226364
rect 186314 226352 186320 226364
rect 148376 226324 186320 226352
rect 148376 226312 148382 226324
rect 186314 226312 186320 226324
rect 186372 226312 186378 226364
rect 157978 225020 157984 225072
rect 158036 225060 158042 225072
rect 186406 225060 186412 225072
rect 158036 225032 186412 225060
rect 158036 225020 158042 225032
rect 186406 225020 186412 225032
rect 186464 225020 186470 225072
rect 133230 224952 133236 225004
rect 133288 224992 133294 225004
rect 186314 224992 186320 225004
rect 133288 224964 186320 224992
rect 133288 224952 133294 224964
rect 186314 224952 186320 224964
rect 186372 224952 186378 225004
rect 151078 223592 151084 223644
rect 151136 223632 151142 223644
rect 186314 223632 186320 223644
rect 151136 223604 186320 223632
rect 151136 223592 151142 223604
rect 186314 223592 186320 223604
rect 186372 223592 186378 223644
rect 145558 222164 145564 222216
rect 145616 222204 145622 222216
rect 186314 222204 186320 222216
rect 145616 222176 186320 222204
rect 145616 222164 145622 222176
rect 186314 222164 186320 222176
rect 186372 222164 186378 222216
rect 162118 220804 162124 220856
rect 162176 220844 162182 220856
rect 186314 220844 186320 220856
rect 162176 220816 186320 220844
rect 162176 220804 162182 220816
rect 186314 220804 186320 220816
rect 186372 220804 186378 220856
rect 145650 219444 145656 219496
rect 145708 219484 145714 219496
rect 186314 219484 186320 219496
rect 145708 219456 186320 219484
rect 145708 219444 145714 219456
rect 186314 219444 186320 219456
rect 186372 219444 186378 219496
rect 156598 218084 156604 218136
rect 156656 218124 156662 218136
rect 186406 218124 186412 218136
rect 156656 218096 186412 218124
rect 156656 218084 156662 218096
rect 186406 218084 186412 218096
rect 186464 218084 186470 218136
rect 135898 218016 135904 218068
rect 135956 218056 135962 218068
rect 186314 218056 186320 218068
rect 135956 218028 186320 218056
rect 135956 218016 135962 218028
rect 186314 218016 186320 218028
rect 186372 218016 186378 218068
rect 542998 218016 543004 218068
rect 543056 218056 543062 218068
rect 580166 218056 580172 218068
rect 543056 218028 580172 218056
rect 543056 218016 543062 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 149698 216656 149704 216708
rect 149756 216696 149762 216708
rect 186314 216696 186320 216708
rect 149756 216668 186320 216696
rect 149756 216656 149762 216668
rect 186314 216656 186320 216668
rect 186372 216656 186378 216708
rect 142798 215296 142804 215348
rect 142856 215336 142862 215348
rect 186314 215336 186320 215348
rect 142856 215308 186320 215336
rect 142856 215296 142862 215308
rect 186314 215296 186320 215308
rect 186372 215296 186378 215348
rect 155218 213936 155224 213988
rect 155276 213976 155282 213988
rect 186314 213976 186320 213988
rect 155276 213948 186320 213976
rect 155276 213936 155282 213948
rect 186314 213936 186320 213948
rect 186372 213936 186378 213988
rect 135990 212508 135996 212560
rect 136048 212548 136054 212560
rect 186314 212548 186320 212560
rect 136048 212520 186320 212548
rect 136048 212508 136054 212520
rect 186314 212508 186320 212520
rect 186372 212508 186378 212560
rect 145742 211148 145748 211200
rect 145800 211188 145806 211200
rect 186314 211188 186320 211200
rect 145800 211160 186320 211188
rect 145800 211148 145806 211160
rect 186314 211148 186320 211160
rect 186372 211148 186378 211200
rect 160738 209856 160744 209908
rect 160796 209896 160802 209908
rect 186314 209896 186320 209908
rect 160796 209868 186320 209896
rect 160796 209856 160802 209868
rect 186314 209856 186320 209868
rect 186372 209856 186378 209908
rect 149790 209788 149796 209840
rect 149848 209828 149854 209840
rect 186406 209828 186412 209840
rect 149848 209800 186412 209828
rect 149848 209788 149854 209800
rect 186406 209788 186412 209800
rect 186464 209788 186470 209840
rect 159358 207000 159364 207052
rect 159416 207040 159422 207052
rect 186314 207040 186320 207052
rect 159416 207012 186320 207040
rect 159416 207000 159422 207012
rect 186314 207000 186320 207012
rect 186372 207000 186378 207052
rect 158070 205640 158076 205692
rect 158128 205680 158134 205692
rect 186314 205680 186320 205692
rect 158128 205652 186320 205680
rect 158128 205640 158134 205652
rect 186314 205640 186320 205652
rect 186372 205640 186378 205692
rect 140038 204280 140044 204332
rect 140096 204320 140102 204332
rect 186314 204320 186320 204332
rect 140096 204292 186320 204320
rect 140096 204280 140102 204292
rect 186314 204280 186320 204292
rect 186372 204280 186378 204332
rect 146938 202920 146944 202972
rect 146996 202960 147002 202972
rect 186314 202960 186320 202972
rect 146996 202932 186320 202960
rect 146996 202920 147002 202932
rect 186314 202920 186320 202932
rect 186372 202920 186378 202972
rect 134610 202852 134616 202904
rect 134668 202892 134674 202904
rect 186406 202892 186412 202904
rect 134668 202864 186412 202892
rect 134668 202852 134674 202864
rect 186406 202852 186412 202864
rect 186464 202852 186470 202904
rect 411254 202852 411260 202904
rect 411312 202892 411318 202904
rect 540238 202892 540244 202904
rect 411312 202864 540244 202892
rect 411312 202852 411318 202864
rect 540238 202852 540244 202864
rect 540296 202852 540302 202904
rect 411254 201560 411260 201612
rect 411312 201600 411318 201612
rect 414658 201600 414664 201612
rect 411312 201572 414664 201600
rect 411312 201560 411318 201572
rect 414658 201560 414664 201572
rect 414716 201560 414722 201612
rect 134518 201492 134524 201544
rect 134576 201532 134582 201544
rect 186314 201532 186320 201544
rect 134576 201504 186320 201532
rect 134576 201492 134582 201504
rect 186314 201492 186320 201504
rect 186372 201492 186378 201544
rect 144178 200132 144184 200184
rect 144236 200172 144242 200184
rect 186314 200172 186320 200184
rect 144236 200144 186320 200172
rect 144236 200132 144242 200144
rect 186314 200132 186320 200144
rect 186372 200132 186378 200184
rect 134702 198704 134708 198756
rect 134760 198744 134766 198756
rect 186314 198744 186320 198756
rect 134760 198716 186320 198744
rect 134760 198704 134766 198716
rect 186314 198704 186320 198716
rect 186372 198704 186378 198756
rect 411254 198704 411260 198756
rect 411312 198744 411318 198756
rect 540330 198744 540336 198756
rect 411312 198716 540336 198744
rect 411312 198704 411318 198716
rect 540330 198704 540336 198716
rect 540388 198704 540394 198756
rect 159450 197344 159456 197396
rect 159508 197384 159514 197396
rect 186314 197384 186320 197396
rect 159508 197356 186320 197384
rect 159508 197344 159514 197356
rect 186314 197344 186320 197356
rect 186372 197344 186378 197396
rect 411254 197344 411260 197396
rect 411312 197384 411318 197396
rect 540422 197384 540428 197396
rect 411312 197356 540428 197384
rect 411312 197344 411318 197356
rect 540422 197344 540428 197356
rect 540480 197344 540486 197396
rect 147030 194624 147036 194676
rect 147088 194664 147094 194676
rect 186314 194664 186320 194676
rect 147088 194636 186320 194664
rect 147088 194624 147094 194636
rect 186314 194624 186320 194636
rect 186372 194624 186378 194676
rect 141418 194556 141424 194608
rect 141476 194596 141482 194608
rect 186406 194596 186412 194608
rect 141476 194568 186412 194596
rect 141476 194556 141482 194568
rect 186406 194556 186412 194568
rect 186464 194556 186470 194608
rect 411254 193536 411260 193588
rect 411312 193576 411318 193588
rect 413370 193576 413376 193588
rect 411312 193548 413376 193576
rect 411312 193536 411318 193548
rect 413370 193536 413376 193548
rect 413428 193536 413434 193588
rect 137278 193196 137284 193248
rect 137336 193236 137342 193248
rect 186314 193236 186320 193248
rect 137336 193208 186320 193236
rect 137336 193196 137342 193208
rect 186314 193196 186320 193208
rect 186372 193196 186378 193248
rect 147122 191836 147128 191888
rect 147180 191876 147186 191888
rect 186314 191876 186320 191888
rect 147180 191848 186320 191876
rect 147180 191836 147186 191848
rect 186314 191836 186320 191848
rect 186372 191836 186378 191888
rect 93670 191224 93676 191276
rect 93728 191264 93734 191276
rect 166258 191264 166264 191276
rect 93728 191236 166264 191264
rect 93728 191224 93734 191236
rect 166258 191224 166264 191236
rect 166316 191224 166322 191276
rect 92382 191156 92388 191208
rect 92440 191196 92446 191208
rect 188338 191196 188344 191208
rect 92440 191168 188344 191196
rect 92440 191156 92446 191168
rect 188338 191156 188344 191168
rect 188396 191156 188402 191208
rect 79962 191088 79968 191140
rect 80020 191128 80026 191140
rect 189718 191128 189724 191140
rect 80020 191100 189724 191128
rect 80020 191088 80026 191100
rect 189718 191088 189724 191100
rect 189776 191088 189782 191140
rect 140130 190476 140136 190528
rect 140188 190516 140194 190528
rect 186314 190516 186320 190528
rect 140188 190488 186320 190516
rect 140188 190476 140194 190488
rect 186314 190476 186320 190488
rect 186372 190476 186378 190528
rect 156690 189048 156696 189100
rect 156748 189088 156754 189100
rect 186314 189088 186320 189100
rect 156748 189060 186320 189088
rect 156748 189048 156754 189060
rect 186314 189048 186320 189060
rect 186372 189048 186378 189100
rect 411254 189048 411260 189100
rect 411312 189088 411318 189100
rect 428458 189088 428464 189100
rect 411312 189060 428464 189088
rect 411312 189048 411318 189060
rect 428458 189048 428464 189060
rect 428516 189048 428522 189100
rect 159542 187756 159548 187808
rect 159600 187796 159606 187808
rect 186406 187796 186412 187808
rect 159600 187768 186412 187796
rect 159600 187756 159606 187768
rect 186406 187756 186412 187768
rect 186464 187756 186470 187808
rect 133322 187688 133328 187740
rect 133380 187728 133386 187740
rect 186314 187728 186320 187740
rect 133380 187700 186320 187728
rect 133380 187688 133386 187700
rect 186314 187688 186320 187700
rect 186372 187688 186378 187740
rect 411254 187688 411260 187740
rect 411312 187728 411318 187740
rect 428550 187728 428556 187740
rect 411312 187700 428556 187728
rect 411312 187688 411318 187700
rect 428550 187688 428556 187700
rect 428608 187688 428614 187740
rect 137370 186328 137376 186380
rect 137428 186368 137434 186380
rect 186314 186368 186320 186380
rect 137428 186340 186320 186368
rect 137428 186328 137434 186340
rect 186314 186328 186320 186340
rect 186372 186328 186378 186380
rect 411254 186328 411260 186380
rect 411312 186368 411318 186380
rect 418982 186368 418988 186380
rect 411312 186340 418988 186368
rect 411312 186328 411318 186340
rect 418982 186328 418988 186340
rect 419040 186328 419046 186380
rect 141510 184900 141516 184952
rect 141568 184940 141574 184952
rect 186314 184940 186320 184952
rect 141568 184912 186320 184940
rect 141568 184900 141574 184912
rect 186314 184900 186320 184912
rect 186372 184900 186378 184952
rect 140222 183540 140228 183592
rect 140280 183580 140286 183592
rect 186314 183580 186320 183592
rect 140280 183552 186320 183580
rect 140280 183540 140286 183552
rect 186314 183540 186320 183552
rect 186372 183540 186378 183592
rect 411254 183540 411260 183592
rect 411312 183580 411318 183592
rect 428642 183580 428648 183592
rect 411312 183552 428648 183580
rect 411312 183540 411318 183552
rect 428642 183540 428648 183552
rect 428700 183540 428706 183592
rect 156874 182180 156880 182232
rect 156932 182220 156938 182232
rect 186314 182220 186320 182232
rect 156932 182192 186320 182220
rect 156932 182180 156938 182192
rect 186314 182180 186320 182192
rect 186372 182180 186378 182232
rect 411254 182180 411260 182232
rect 411312 182220 411318 182232
rect 436738 182220 436744 182232
rect 411312 182192 436744 182220
rect 411312 182180 411318 182192
rect 436738 182180 436744 182192
rect 436796 182180 436802 182232
rect 156782 180888 156788 180940
rect 156840 180928 156846 180940
rect 186314 180928 186320 180940
rect 156840 180900 186320 180928
rect 156840 180888 156846 180900
rect 186314 180888 186320 180900
rect 186372 180888 186378 180940
rect 140314 180820 140320 180872
rect 140372 180860 140378 180872
rect 186406 180860 186412 180872
rect 140372 180832 186412 180860
rect 140372 180820 140378 180832
rect 186406 180820 186412 180832
rect 186464 180820 186470 180872
rect 137462 179392 137468 179444
rect 137520 179432 137526 179444
rect 186314 179432 186320 179444
rect 137520 179404 186320 179432
rect 137520 179392 137526 179404
rect 186314 179392 186320 179404
rect 186372 179392 186378 179444
rect 411254 179392 411260 179444
rect 411312 179432 411318 179444
rect 425698 179432 425704 179444
rect 411312 179404 425704 179432
rect 411312 179392 411318 179404
rect 425698 179392 425704 179404
rect 425756 179392 425762 179444
rect 144270 178032 144276 178084
rect 144328 178072 144334 178084
rect 186314 178072 186320 178084
rect 144328 178044 186320 178072
rect 144328 178032 144334 178044
rect 186314 178032 186320 178044
rect 186372 178032 186378 178084
rect 411254 178032 411260 178084
rect 411312 178072 411318 178084
rect 435358 178072 435364 178084
rect 411312 178044 435364 178072
rect 411312 178032 411318 178044
rect 435358 178032 435364 178044
rect 435416 178032 435422 178084
rect 543090 178032 543096 178084
rect 543148 178072 543154 178084
rect 580166 178072 580172 178084
rect 543148 178044 580172 178072
rect 543148 178032 543154 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 138658 176672 138664 176724
rect 138716 176712 138722 176724
rect 186314 176712 186320 176724
rect 138716 176684 186320 176712
rect 138716 176672 138722 176684
rect 186314 176672 186320 176684
rect 186372 176672 186378 176724
rect 411254 176672 411260 176724
rect 411312 176712 411318 176724
rect 417418 176712 417424 176724
rect 411312 176684 417424 176712
rect 411312 176672 411318 176684
rect 417418 176672 417424 176684
rect 417476 176672 417482 176724
rect 141602 175244 141608 175296
rect 141660 175284 141666 175296
rect 186314 175284 186320 175296
rect 141660 175256 186320 175284
rect 141660 175244 141666 175256
rect 186314 175244 186320 175256
rect 186372 175244 186378 175296
rect 411254 174428 411260 174480
rect 411312 174468 411318 174480
rect 414934 174468 414940 174480
rect 411312 174440 414940 174468
rect 411312 174428 411318 174440
rect 414934 174428 414940 174440
rect 414992 174428 414998 174480
rect 164970 173884 164976 173936
rect 165028 173924 165034 173936
rect 186314 173924 186320 173936
rect 165028 173896 186320 173924
rect 165028 173884 165034 173896
rect 186314 173884 186320 173896
rect 186372 173884 186378 173936
rect 160830 172592 160836 172644
rect 160888 172632 160894 172644
rect 186314 172632 186320 172644
rect 160888 172604 186320 172632
rect 160888 172592 160894 172604
rect 186314 172592 186320 172604
rect 186372 172592 186378 172644
rect 138750 172524 138756 172576
rect 138808 172564 138814 172576
rect 186406 172564 186412 172576
rect 138808 172536 186412 172564
rect 138808 172524 138814 172536
rect 186406 172524 186412 172536
rect 186464 172524 186470 172576
rect 411254 172524 411260 172576
rect 411312 172564 411318 172576
rect 432598 172564 432604 172576
rect 411312 172536 432604 172564
rect 411312 172524 411318 172536
rect 432598 172524 432604 172536
rect 432656 172524 432662 172576
rect 137554 171096 137560 171148
rect 137612 171136 137618 171148
rect 186314 171136 186320 171148
rect 137612 171108 186320 171136
rect 137612 171096 137618 171108
rect 186314 171096 186320 171108
rect 186372 171096 186378 171148
rect 411254 171096 411260 171148
rect 411312 171136 411318 171148
rect 431218 171136 431224 171148
rect 411312 171108 431224 171136
rect 411312 171096 411318 171108
rect 431218 171096 431224 171108
rect 431276 171096 431282 171148
rect 131850 169736 131856 169788
rect 131908 169776 131914 169788
rect 186314 169776 186320 169788
rect 131908 169748 186320 169776
rect 131908 169736 131914 169748
rect 186314 169736 186320 169748
rect 186372 169736 186378 169788
rect 158162 168376 158168 168428
rect 158220 168416 158226 168428
rect 186314 168416 186320 168428
rect 158220 168388 186320 168416
rect 158220 168376 158226 168388
rect 186314 168376 186320 168388
rect 186372 168376 186378 168428
rect 411254 168376 411260 168428
rect 411312 168416 411318 168428
rect 429838 168416 429844 168428
rect 411312 168388 429844 168416
rect 411312 168376 411318 168388
rect 429838 168376 429844 168388
rect 429896 168376 429902 168428
rect 162210 167016 162216 167068
rect 162268 167056 162274 167068
rect 186314 167056 186320 167068
rect 162268 167028 186320 167056
rect 162268 167016 162274 167028
rect 186314 167016 186320 167028
rect 186372 167016 186378 167068
rect 411254 167016 411260 167068
rect 411312 167056 411318 167068
rect 428734 167056 428740 167068
rect 411312 167028 428740 167056
rect 411312 167016 411318 167028
rect 428734 167016 428740 167028
rect 428792 167016 428798 167068
rect 159634 165656 159640 165708
rect 159692 165696 159698 165708
rect 186314 165696 186320 165708
rect 159692 165668 186320 165696
rect 159692 165656 159698 165668
rect 186314 165656 186320 165668
rect 186372 165656 186378 165708
rect 158254 165588 158260 165640
rect 158312 165628 158318 165640
rect 186406 165628 186412 165640
rect 158312 165600 186412 165628
rect 158312 165588 158318 165600
rect 186406 165588 186412 165600
rect 186464 165588 186470 165640
rect 155310 164228 155316 164280
rect 155368 164268 155374 164280
rect 186314 164268 186320 164280
rect 155368 164240 186320 164268
rect 155368 164228 155374 164240
rect 186314 164228 186320 164240
rect 186372 164228 186378 164280
rect 411254 164228 411260 164280
rect 411312 164268 411318 164280
rect 425790 164268 425796 164280
rect 411312 164240 425796 164268
rect 411312 164228 411318 164240
rect 425790 164228 425796 164240
rect 425848 164228 425854 164280
rect 160922 162868 160928 162920
rect 160980 162908 160986 162920
rect 186314 162908 186320 162920
rect 160980 162880 186320 162908
rect 160980 162868 160986 162880
rect 186314 162868 186320 162880
rect 186372 162868 186378 162920
rect 411254 162868 411260 162920
rect 411312 162908 411318 162920
rect 424318 162908 424324 162920
rect 411312 162880 424324 162908
rect 411312 162868 411318 162880
rect 424318 162868 424324 162880
rect 424376 162868 424382 162920
rect 134794 161440 134800 161492
rect 134852 161480 134858 161492
rect 186314 161480 186320 161492
rect 134852 161452 186320 161480
rect 134852 161440 134858 161452
rect 186314 161440 186320 161452
rect 186372 161440 186378 161492
rect 411254 161440 411260 161492
rect 411312 161480 411318 161492
rect 424410 161480 424416 161492
rect 411312 161452 424416 161480
rect 411312 161440 411318 161452
rect 424410 161440 424416 161452
rect 424468 161440 424474 161492
rect 158346 160080 158352 160132
rect 158404 160120 158410 160132
rect 186314 160120 186320 160132
rect 158404 160092 186320 160120
rect 158404 160080 158410 160092
rect 186314 160080 186320 160092
rect 186372 160080 186378 160132
rect 133506 158720 133512 158772
rect 133564 158760 133570 158772
rect 186314 158760 186320 158772
rect 133564 158732 186320 158760
rect 133564 158720 133570 158732
rect 186314 158720 186320 158732
rect 186372 158720 186378 158772
rect 411254 158720 411260 158772
rect 411312 158760 411318 158772
rect 423122 158760 423128 158772
rect 411312 158732 423128 158760
rect 411312 158720 411318 158732
rect 423122 158720 423128 158732
rect 423180 158720 423186 158772
rect 156966 157428 156972 157480
rect 157024 157468 157030 157480
rect 186406 157468 186412 157480
rect 157024 157440 186412 157468
rect 157024 157428 157030 157440
rect 186406 157428 186412 157440
rect 186464 157428 186470 157480
rect 133414 157360 133420 157412
rect 133472 157400 133478 157412
rect 186314 157400 186320 157412
rect 133472 157372 186320 157400
rect 133472 157360 133478 157372
rect 186314 157360 186320 157372
rect 186372 157360 186378 157412
rect 411254 157360 411260 157412
rect 411312 157400 411318 157412
rect 425882 157400 425888 157412
rect 411312 157372 425888 157400
rect 411312 157360 411318 157372
rect 425882 157360 425888 157372
rect 425940 157360 425946 157412
rect 136082 155932 136088 155984
rect 136140 155972 136146 155984
rect 186314 155972 186320 155984
rect 136140 155944 186320 155972
rect 136140 155932 136146 155944
rect 186314 155932 186320 155944
rect 186372 155932 186378 155984
rect 411254 155932 411260 155984
rect 411312 155972 411318 155984
rect 423030 155972 423036 155984
rect 411312 155944 423036 155972
rect 411312 155932 411318 155944
rect 423030 155932 423036 155944
rect 423088 155932 423094 155984
rect 133598 154572 133604 154624
rect 133656 154612 133662 154624
rect 186314 154612 186320 154624
rect 133656 154584 186320 154612
rect 133656 154572 133662 154584
rect 186314 154572 186320 154584
rect 186372 154572 186378 154624
rect 138842 153212 138848 153264
rect 138900 153252 138906 153264
rect 186314 153252 186320 153264
rect 138900 153224 186320 153252
rect 138900 153212 138906 153224
rect 186314 153212 186320 153224
rect 186372 153212 186378 153264
rect 411254 153212 411260 153264
rect 411312 153252 411318 153264
rect 417510 153252 417516 153264
rect 411312 153224 417516 153252
rect 411312 153212 411318 153224
rect 417510 153212 417516 153224
rect 417568 153212 417574 153264
rect 141694 151784 141700 151836
rect 141752 151824 141758 151836
rect 186314 151824 186320 151836
rect 141752 151796 186320 151824
rect 141752 151784 141758 151796
rect 186314 151784 186320 151796
rect 186372 151784 186378 151836
rect 411254 151784 411260 151836
rect 411312 151824 411318 151836
rect 422938 151824 422944 151836
rect 411312 151796 422944 151824
rect 411312 151784 411318 151796
rect 422938 151784 422944 151796
rect 422996 151784 423002 151836
rect 166350 150492 166356 150544
rect 166408 150532 166414 150544
rect 186406 150532 186412 150544
rect 166408 150504 186412 150532
rect 166408 150492 166414 150504
rect 186406 150492 186412 150504
rect 186464 150492 186470 150544
rect 155402 150424 155408 150476
rect 155460 150464 155466 150476
rect 186314 150464 186320 150476
rect 155460 150436 186320 150464
rect 155460 150424 155466 150436
rect 186314 150424 186320 150436
rect 186372 150424 186378 150476
rect 151170 149064 151176 149116
rect 151228 149104 151234 149116
rect 186314 149104 186320 149116
rect 151228 149076 186320 149104
rect 151228 149064 151234 149076
rect 186314 149064 186320 149076
rect 186372 149064 186378 149116
rect 411254 149064 411260 149116
rect 411312 149104 411318 149116
rect 417602 149104 417608 149116
rect 411312 149076 417608 149104
rect 411312 149064 411318 149076
rect 417602 149064 417608 149076
rect 417660 149064 417666 149116
rect 144362 147636 144368 147688
rect 144420 147676 144426 147688
rect 186314 147676 186320 147688
rect 144420 147648 186320 147676
rect 144420 147636 144426 147648
rect 186314 147636 186320 147648
rect 186372 147636 186378 147688
rect 411254 147636 411260 147688
rect 411312 147676 411318 147688
rect 421650 147676 421656 147688
rect 411312 147648 421656 147676
rect 411312 147636 411318 147648
rect 421650 147636 421656 147648
rect 421708 147636 421714 147688
rect 155494 146276 155500 146328
rect 155552 146316 155558 146328
rect 186314 146316 186320 146328
rect 155552 146288 186320 146316
rect 155552 146276 155558 146288
rect 186314 146276 186320 146288
rect 186372 146276 186378 146328
rect 411254 146276 411260 146328
rect 411312 146316 411318 146328
rect 419166 146316 419172 146328
rect 411312 146288 419172 146316
rect 411312 146276 411318 146288
rect 419166 146276 419172 146288
rect 419224 146276 419230 146328
rect 151262 144916 151268 144968
rect 151320 144956 151326 144968
rect 186314 144956 186320 144968
rect 151320 144928 186320 144956
rect 151320 144916 151326 144928
rect 186314 144916 186320 144928
rect 186372 144916 186378 144968
rect 152458 143624 152464 143676
rect 152516 143664 152522 143676
rect 186314 143664 186320 143676
rect 152516 143636 186320 143664
rect 152516 143624 152522 143636
rect 186314 143624 186320 143636
rect 186372 143624 186378 143676
rect 144454 143556 144460 143608
rect 144512 143596 144518 143608
rect 186406 143596 186412 143608
rect 144512 143568 186412 143596
rect 144512 143556 144518 143568
rect 186406 143556 186412 143568
rect 186464 143556 186470 143608
rect 411254 143556 411260 143608
rect 411312 143596 411318 143608
rect 421558 143596 421564 143608
rect 411312 143568 421564 143596
rect 411312 143556 411318 143568
rect 421558 143556 421564 143568
rect 421616 143556 421622 143608
rect 148410 142128 148416 142180
rect 148468 142168 148474 142180
rect 186314 142168 186320 142180
rect 148468 142140 186320 142168
rect 148468 142128 148474 142140
rect 186314 142128 186320 142140
rect 186372 142128 186378 142180
rect 411254 142128 411260 142180
rect 411312 142168 411318 142180
rect 429930 142168 429936 142180
rect 411312 142140 429936 142168
rect 411312 142128 411318 142140
rect 429930 142128 429936 142140
rect 429988 142128 429994 142180
rect 411254 140768 411260 140820
rect 411312 140808 411318 140820
rect 417694 140808 417700 140820
rect 411312 140780 417700 140808
rect 411312 140768 411318 140780
rect 417694 140768 417700 140780
rect 417752 140768 417758 140820
rect 152550 139408 152556 139460
rect 152608 139448 152614 139460
rect 186314 139448 186320 139460
rect 152608 139420 186320 139448
rect 152608 139408 152614 139420
rect 186314 139408 186320 139420
rect 186372 139408 186378 139460
rect 414658 139340 414664 139392
rect 414716 139380 414722 139392
rect 580166 139380 580172 139392
rect 414716 139352 580172 139380
rect 414716 139340 414722 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 148502 137980 148508 138032
rect 148560 138020 148566 138032
rect 186314 138020 186320 138032
rect 148560 137992 186320 138020
rect 148560 137980 148566 137992
rect 186314 137980 186320 137992
rect 186372 137980 186378 138032
rect 411254 137980 411260 138032
rect 411312 138020 411318 138032
rect 426066 138020 426072 138032
rect 411312 137992 426072 138020
rect 411312 137980 411318 137992
rect 426066 137980 426072 137992
rect 426124 137980 426130 138032
rect 142890 136620 142896 136672
rect 142948 136660 142954 136672
rect 186314 136660 186320 136672
rect 142948 136632 186320 136660
rect 142948 136620 142954 136632
rect 186314 136620 186320 136632
rect 186372 136620 186378 136672
rect 411254 136620 411260 136672
rect 411312 136660 411318 136672
rect 425974 136660 425980 136672
rect 411312 136632 425980 136660
rect 411312 136620 411318 136632
rect 425974 136620 425980 136632
rect 426032 136620 426038 136672
rect 152642 135328 152648 135380
rect 152700 135368 152706 135380
rect 186406 135368 186412 135380
rect 152700 135340 186412 135368
rect 152700 135328 152706 135340
rect 186406 135328 186412 135340
rect 186464 135328 186470 135380
rect 148594 135260 148600 135312
rect 148652 135300 148658 135312
rect 186314 135300 186320 135312
rect 148652 135272 186320 135300
rect 148652 135260 148658 135272
rect 186314 135260 186320 135272
rect 186372 135260 186378 135312
rect 411254 135260 411260 135312
rect 411312 135300 411318 135312
rect 431310 135300 431316 135312
rect 411312 135272 431316 135300
rect 411312 135260 411318 135272
rect 431310 135260 431316 135272
rect 431368 135260 431374 135312
rect 93762 133288 93768 133340
rect 93820 133328 93826 133340
rect 164878 133328 164884 133340
rect 93820 133300 164884 133328
rect 93820 133288 93826 133300
rect 164878 133288 164884 133300
rect 164936 133288 164942 133340
rect 117222 133220 117228 133272
rect 117280 133260 117286 133272
rect 188522 133260 188528 133272
rect 117280 133232 188528 133260
rect 117280 133220 117286 133232
rect 188522 133220 188528 133232
rect 188580 133220 188586 133272
rect 113082 133152 113088 133204
rect 113140 133192 113146 133204
rect 188430 133192 188436 133204
rect 113140 133164 188436 133192
rect 113140 133152 113146 133164
rect 188430 133152 188436 133164
rect 188488 133152 188494 133204
rect 152734 132472 152740 132524
rect 152792 132512 152798 132524
rect 186314 132512 186320 132524
rect 152792 132484 186320 132512
rect 152792 132472 152798 132484
rect 186314 132472 186320 132484
rect 186372 132472 186378 132524
rect 411254 132472 411260 132524
rect 411312 132512 411318 132524
rect 424502 132512 424508 132524
rect 411312 132484 424508 132512
rect 411312 132472 411318 132484
rect 424502 132472 424508 132484
rect 424560 132472 424566 132524
rect 110322 131860 110328 131912
rect 110380 131900 110386 131912
rect 189994 131900 190000 131912
rect 110380 131872 190000 131900
rect 110380 131860 110386 131872
rect 189994 131860 190000 131872
rect 190052 131860 190058 131912
rect 97902 131792 97908 131844
rect 97960 131832 97966 131844
rect 189902 131832 189908 131844
rect 97960 131804 189908 131832
rect 97960 131792 97966 131804
rect 189902 131792 189908 131804
rect 189960 131792 189966 131844
rect 48130 131724 48136 131776
rect 48188 131764 48194 131776
rect 189810 131764 189816 131776
rect 48188 131736 189816 131764
rect 48188 131724 48194 131736
rect 189810 131724 189816 131736
rect 189868 131724 189874 131776
rect 413462 131452 413468 131504
rect 413520 131492 413526 131504
rect 521746 131492 521752 131504
rect 413520 131464 521752 131492
rect 413520 131452 413526 131464
rect 521746 131452 521752 131464
rect 521804 131452 521810 131504
rect 439682 131384 439688 131436
rect 439740 131424 439746 131436
rect 472066 131424 472072 131436
rect 439740 131396 472072 131424
rect 439740 131384 439746 131396
rect 472066 131384 472072 131396
rect 472124 131384 472130 131436
rect 414658 131316 414664 131368
rect 414716 131356 414722 131368
rect 478874 131356 478880 131368
rect 414716 131328 478880 131356
rect 414716 131316 414722 131328
rect 478874 131316 478880 131328
rect 478932 131316 478938 131368
rect 414750 131248 414756 131300
rect 414808 131288 414814 131300
rect 485958 131288 485964 131300
rect 414808 131260 485964 131288
rect 414808 131248 414814 131260
rect 485958 131248 485964 131260
rect 486016 131248 486022 131300
rect 1302 131180 1308 131232
rect 1360 131220 1366 131232
rect 55122 131220 55128 131232
rect 1360 131192 55128 131220
rect 1360 131180 1366 131192
rect 55122 131180 55128 131192
rect 55180 131180 55186 131232
rect 438118 131180 438124 131232
rect 438176 131220 438182 131232
rect 536006 131220 536012 131232
rect 438176 131192 536012 131220
rect 438176 131180 438182 131192
rect 536006 131180 536012 131192
rect 536064 131180 536070 131232
rect 2682 131112 2688 131164
rect 2740 131152 2746 131164
rect 104894 131152 104900 131164
rect 2740 131124 104900 131152
rect 2740 131112 2746 131124
rect 104894 131112 104900 131124
rect 104952 131112 104958 131164
rect 148686 131112 148692 131164
rect 148744 131152 148750 131164
rect 186314 131152 186320 131164
rect 148744 131124 186320 131152
rect 148744 131112 148750 131124
rect 186314 131112 186320 131124
rect 186372 131112 186378 131164
rect 411254 131112 411260 131164
rect 411312 131152 411318 131164
rect 415026 131152 415032 131164
rect 411312 131124 415032 131152
rect 411312 131112 411318 131124
rect 415026 131112 415032 131124
rect 415084 131112 415090 131164
rect 439498 131112 439504 131164
rect 439556 131152 439562 131164
rect 443178 131152 443184 131164
rect 439556 131124 443184 131152
rect 439556 131112 439562 131124
rect 443178 131112 443184 131124
rect 443236 131112 443242 131164
rect 48038 130500 48044 130552
rect 48096 130540 48102 130552
rect 133138 130540 133144 130552
rect 48096 130512 133144 130540
rect 48096 130500 48102 130512
rect 133138 130500 133144 130512
rect 133196 130500 133202 130552
rect 78582 130432 78588 130484
rect 78640 130472 78646 130484
rect 190178 130472 190184 130484
rect 78640 130444 190184 130472
rect 78640 130432 78646 130444
rect 190178 130432 190184 130444
rect 190236 130432 190242 130484
rect 439866 130432 439872 130484
rect 439924 130472 439930 130484
rect 542538 130472 542544 130484
rect 439924 130444 542544 130472
rect 439924 130432 439930 130444
rect 542538 130432 542544 130444
rect 542596 130432 542602 130484
rect 48222 130364 48228 130416
rect 48280 130404 48286 130416
rect 190086 130404 190092 130416
rect 48280 130376 190092 130404
rect 48280 130364 48286 130376
rect 190086 130364 190092 130376
rect 190144 130364 190150 130416
rect 438762 130364 438768 130416
rect 438820 130404 438826 130416
rect 450262 130404 450268 130416
rect 438820 130376 450268 130404
rect 438820 130364 438826 130376
rect 450262 130364 450268 130376
rect 450320 130364 450326 130416
rect 439590 130296 439596 130348
rect 439648 130336 439654 130348
rect 464522 130336 464528 130348
rect 439648 130308 464528 130336
rect 439648 130296 439654 130308
rect 464522 130296 464528 130308
rect 464580 130296 464586 130348
rect 419074 130228 419080 130280
rect 419132 130268 419138 130280
rect 493134 130268 493140 130280
rect 419132 130240 493140 130268
rect 419132 130228 419138 130240
rect 493134 130228 493140 130240
rect 493192 130228 493198 130280
rect 439774 130160 439780 130212
rect 439832 130200 439838 130212
rect 514892 130200 514898 130212
rect 439832 130172 514898 130200
rect 439832 130160 439838 130172
rect 514892 130160 514898 130172
rect 514950 130160 514956 130212
rect 420178 130092 420184 130144
rect 420236 130132 420242 130144
rect 500632 130132 500638 130144
rect 420236 130104 500638 130132
rect 420236 130092 420242 130104
rect 500632 130092 500638 130104
rect 500690 130092 500696 130144
rect 420270 130024 420276 130076
rect 420328 130064 420334 130076
rect 507394 130064 507400 130076
rect 420328 130036 507400 130064
rect 420328 130024 420334 130036
rect 507394 130024 507400 130036
rect 507452 130024 507458 130076
rect 435542 129956 435548 130008
rect 435600 129996 435606 130008
rect 528830 129996 528836 130008
rect 435600 129968 528836 129996
rect 435600 129956 435606 129968
rect 528830 129956 528836 129968
rect 528888 129956 528894 130008
rect 439958 129888 439964 129940
rect 440016 129928 440022 129940
rect 539318 129928 539324 129940
rect 440016 129900 539324 129928
rect 440016 129888 440022 129900
rect 539318 129888 539324 129900
rect 539376 129888 539382 129940
rect 418798 129820 418804 129872
rect 418856 129860 418862 129872
rect 457438 129860 457444 129872
rect 418856 129832 457444 129860
rect 418856 129820 418862 129832
rect 457438 129820 457444 129832
rect 457496 129820 457502 129872
rect 142982 129752 142988 129804
rect 143040 129792 143046 129804
rect 186314 129792 186320 129804
rect 143040 129764 186320 129792
rect 143040 129752 143046 129764
rect 186314 129752 186320 129764
rect 186372 129752 186378 129804
rect 412266 129752 412272 129804
rect 412324 129792 412330 129804
rect 542354 129792 542360 129804
rect 412324 129764 542360 129792
rect 412324 129752 412330 129764
rect 542354 129752 542360 129764
rect 542412 129752 542418 129804
rect 131114 129684 131120 129736
rect 131172 129724 131178 129736
rect 169018 129724 169024 129736
rect 131172 129696 169024 129724
rect 131172 129684 131178 129696
rect 169018 129684 169024 129696
rect 169076 129684 169082 129736
rect 131298 129616 131304 129668
rect 131356 129656 131362 129668
rect 157978 129656 157984 129668
rect 131356 129628 157984 129656
rect 131356 129616 131362 129628
rect 157978 129616 157984 129628
rect 158036 129616 158042 129668
rect 131206 129548 131212 129600
rect 131264 129588 131270 129600
rect 148318 129588 148324 129600
rect 131264 129560 148324 129588
rect 131264 129548 131270 129560
rect 148318 129548 148324 129560
rect 148376 129548 148382 129600
rect 411254 128460 411260 128512
rect 411312 128500 411318 128512
rect 424594 128500 424600 128512
rect 411312 128472 424600 128500
rect 411312 128460 411318 128472
rect 424594 128460 424600 128472
rect 424652 128460 424658 128512
rect 151354 128392 151360 128444
rect 151412 128432 151418 128444
rect 186406 128432 186412 128444
rect 151412 128404 186412 128432
rect 151412 128392 151418 128404
rect 186406 128392 186412 128404
rect 186464 128392 186470 128444
rect 421926 128392 421932 128444
rect 421984 128432 421990 128444
rect 437474 128432 437480 128444
rect 421984 128404 437480 128432
rect 421984 128392 421990 128404
rect 437474 128392 437480 128404
rect 437532 128392 437538 128444
rect 147214 128324 147220 128376
rect 147272 128364 147278 128376
rect 186314 128364 186320 128376
rect 147272 128336 186320 128364
rect 147272 128324 147278 128336
rect 186314 128324 186320 128336
rect 186372 128324 186378 128376
rect 412358 128324 412364 128376
rect 412416 128364 412422 128376
rect 542446 128364 542452 128376
rect 412416 128336 542452 128364
rect 412416 128324 412422 128336
rect 542446 128324 542452 128336
rect 542504 128324 542510 128376
rect 132034 128256 132040 128308
rect 132092 128296 132098 128308
rect 151078 128296 151084 128308
rect 132092 128268 151084 128296
rect 132092 128256 132098 128268
rect 151078 128256 151084 128268
rect 151136 128256 151142 128308
rect 132218 128188 132224 128240
rect 132276 128228 132282 128240
rect 133230 128228 133236 128240
rect 132276 128200 133236 128228
rect 132276 128188 132282 128200
rect 133230 128188 133236 128200
rect 133288 128188 133294 128240
rect 411254 127032 411260 127084
rect 411312 127072 411318 127084
rect 432690 127072 432696 127084
rect 411312 127044 432696 127072
rect 411312 127032 411318 127044
rect 432690 127032 432696 127044
rect 432748 127032 432754 127084
rect 143074 126964 143080 127016
rect 143132 127004 143138 127016
rect 186314 127004 186320 127016
rect 143132 126976 186320 127004
rect 143132 126964 143138 126976
rect 186314 126964 186320 126976
rect 186372 126964 186378 127016
rect 413554 126964 413560 127016
rect 413612 127004 413618 127016
rect 437474 127004 437480 127016
rect 413612 126976 437480 127004
rect 413612 126964 413618 126976
rect 437474 126964 437480 126976
rect 437532 126964 437538 127016
rect 131114 126896 131120 126948
rect 131172 126936 131178 126948
rect 162118 126936 162124 126948
rect 131172 126908 162124 126936
rect 131172 126896 131178 126908
rect 162118 126896 162124 126908
rect 162176 126896 162182 126948
rect 132034 126828 132040 126880
rect 132092 126868 132098 126880
rect 145650 126868 145656 126880
rect 132092 126840 145656 126868
rect 132092 126828 132098 126840
rect 145650 126828 145656 126840
rect 145708 126828 145714 126880
rect 131206 126760 131212 126812
rect 131264 126800 131270 126812
rect 145558 126800 145564 126812
rect 131264 126772 145564 126800
rect 131264 126760 131270 126772
rect 145558 126760 145564 126772
rect 145616 126760 145622 126812
rect 411254 125672 411260 125724
rect 411312 125712 411318 125724
rect 416038 125712 416044 125724
rect 411312 125684 416044 125712
rect 411312 125672 411318 125684
rect 416038 125672 416044 125684
rect 416096 125672 416102 125724
rect 151078 125604 151084 125656
rect 151136 125644 151142 125656
rect 186314 125644 186320 125656
rect 151136 125616 186320 125644
rect 151136 125604 151142 125616
rect 186314 125604 186320 125616
rect 186372 125604 186378 125656
rect 413646 125604 413652 125656
rect 413704 125644 413710 125656
rect 437474 125644 437480 125656
rect 413704 125616 437480 125644
rect 413704 125604 413710 125616
rect 437474 125604 437480 125616
rect 437532 125604 437538 125656
rect 541618 125604 541624 125656
rect 541676 125644 541682 125656
rect 580166 125644 580172 125656
rect 541676 125616 580172 125644
rect 541676 125604 541682 125616
rect 580166 125604 580172 125616
rect 580224 125604 580230 125656
rect 131114 125536 131120 125588
rect 131172 125576 131178 125588
rect 156598 125576 156604 125588
rect 131172 125548 156604 125576
rect 131172 125536 131178 125548
rect 156598 125536 156604 125548
rect 156656 125536 156662 125588
rect 131206 125468 131212 125520
rect 131264 125508 131270 125520
rect 135898 125508 135904 125520
rect 131264 125480 135904 125508
rect 131264 125468 131270 125480
rect 135898 125468 135904 125480
rect 135956 125468 135962 125520
rect 436094 124448 436100 124500
rect 436152 124488 436158 124500
rect 438762 124488 438768 124500
rect 436152 124460 438768 124488
rect 436152 124448 436158 124460
rect 438762 124448 438768 124460
rect 438820 124448 438826 124500
rect 145558 124176 145564 124228
rect 145616 124216 145622 124228
rect 186314 124216 186320 124228
rect 145616 124188 186320 124216
rect 145616 124176 145622 124188
rect 186314 124176 186320 124188
rect 186372 124176 186378 124228
rect 414842 124176 414848 124228
rect 414900 124216 414906 124228
rect 437474 124216 437480 124228
rect 414900 124188 437480 124216
rect 414900 124176 414906 124188
rect 437474 124176 437480 124188
rect 437532 124176 437538 124228
rect 132218 124108 132224 124160
rect 132276 124148 132282 124160
rect 149698 124148 149704 124160
rect 132276 124120 149704 124148
rect 132276 124108 132282 124120
rect 149698 124108 149704 124120
rect 149756 124108 149762 124160
rect 131114 124040 131120 124092
rect 131172 124080 131178 124092
rect 142798 124080 142804 124092
rect 131172 124052 142804 124080
rect 131172 124040 131178 124052
rect 142798 124040 142804 124052
rect 142856 124040 142862 124092
rect 411254 122816 411260 122868
rect 411312 122856 411318 122868
rect 435450 122856 435456 122868
rect 411312 122828 435456 122856
rect 411312 122816 411318 122828
rect 435450 122816 435456 122828
rect 435508 122816 435514 122868
rect 131206 122748 131212 122800
rect 131264 122788 131270 122800
rect 155218 122788 155224 122800
rect 131264 122760 155224 122788
rect 131264 122748 131270 122760
rect 155218 122748 155224 122760
rect 155276 122748 155282 122800
rect 131114 122680 131120 122732
rect 131172 122720 131178 122732
rect 145742 122720 145748 122732
rect 131172 122692 145748 122720
rect 131172 122680 131178 122692
rect 145742 122680 145748 122692
rect 145800 122680 145806 122732
rect 131206 122612 131212 122664
rect 131264 122652 131270 122664
rect 135990 122652 135996 122664
rect 131264 122624 135996 122652
rect 131264 122612 131270 122624
rect 135990 122612 135996 122624
rect 136048 122612 136054 122664
rect 411254 121524 411260 121576
rect 411312 121564 411318 121576
rect 416130 121564 416136 121576
rect 411312 121536 416136 121564
rect 411312 121524 411318 121536
rect 416130 121524 416136 121536
rect 416188 121524 416194 121576
rect 149698 121456 149704 121508
rect 149756 121496 149762 121508
rect 186314 121496 186320 121508
rect 149756 121468 186320 121496
rect 149756 121456 149762 121468
rect 186314 121456 186320 121468
rect 186372 121456 186378 121508
rect 413278 121456 413284 121508
rect 413336 121496 413342 121508
rect 437474 121496 437480 121508
rect 413336 121468 437480 121496
rect 413336 121456 413342 121468
rect 437474 121456 437480 121468
rect 437532 121456 437538 121508
rect 131942 121388 131948 121440
rect 132000 121428 132006 121440
rect 160738 121428 160744 121440
rect 132000 121400 160744 121428
rect 132000 121388 132006 121400
rect 160738 121388 160744 121400
rect 160796 121388 160802 121440
rect 131206 121320 131212 121372
rect 131264 121360 131270 121372
rect 149790 121360 149796 121372
rect 131264 121332 149796 121360
rect 131264 121320 131270 121332
rect 149790 121320 149796 121332
rect 149848 121320 149854 121372
rect 145742 120164 145748 120216
rect 145800 120204 145806 120216
rect 186406 120204 186412 120216
rect 145800 120176 186412 120204
rect 145800 120164 145806 120176
rect 186406 120164 186412 120176
rect 186464 120164 186470 120216
rect 434070 120164 434076 120216
rect 434128 120204 434134 120216
rect 436002 120204 436008 120216
rect 434128 120176 436008 120204
rect 434128 120164 434134 120176
rect 436002 120164 436008 120176
rect 436060 120164 436066 120216
rect 142798 120096 142804 120148
rect 142856 120136 142862 120148
rect 186314 120136 186320 120148
rect 142856 120108 186320 120136
rect 142856 120096 142862 120108
rect 186314 120096 186320 120108
rect 186372 120096 186378 120148
rect 418890 120096 418896 120148
rect 418948 120136 418954 120148
rect 437474 120136 437480 120148
rect 418948 120108 437480 120136
rect 418948 120096 418954 120108
rect 437474 120096 437480 120108
rect 437532 120096 437538 120148
rect 132218 120028 132224 120080
rect 132276 120068 132282 120080
rect 186958 120068 186964 120080
rect 132276 120040 186964 120068
rect 132276 120028 132282 120040
rect 186958 120028 186964 120040
rect 187016 120028 187022 120080
rect 411990 120028 411996 120080
rect 412048 120068 412054 120080
rect 437566 120068 437572 120080
rect 412048 120040 437572 120068
rect 412048 120028 412054 120040
rect 437566 120028 437572 120040
rect 437624 120028 437630 120080
rect 131114 119960 131120 120012
rect 131172 120000 131178 120012
rect 159358 120000 159364 120012
rect 131172 119972 159364 120000
rect 131172 119960 131178 119972
rect 159358 119960 159364 119972
rect 159416 119960 159422 120012
rect 135898 118668 135904 118720
rect 135956 118708 135962 118720
rect 186314 118708 186320 118720
rect 135956 118680 186320 118708
rect 135956 118668 135962 118680
rect 186314 118668 186320 118680
rect 186372 118668 186378 118720
rect 411254 118668 411260 118720
rect 411312 118708 411318 118720
rect 424686 118708 424692 118720
rect 411312 118680 424692 118708
rect 411312 118668 411318 118680
rect 424686 118668 424692 118680
rect 424744 118668 424750 118720
rect 131206 118600 131212 118652
rect 131264 118640 131270 118652
rect 158070 118640 158076 118652
rect 131264 118612 158076 118640
rect 131264 118600 131270 118612
rect 158070 118600 158076 118612
rect 158128 118600 158134 118652
rect 413370 118600 413376 118652
rect 413428 118640 413434 118652
rect 437474 118640 437480 118652
rect 413428 118612 437480 118640
rect 413428 118600 413434 118612
rect 437474 118600 437480 118612
rect 437532 118600 437538 118652
rect 131114 118532 131120 118584
rect 131172 118572 131178 118584
rect 140038 118572 140044 118584
rect 131172 118544 140044 118572
rect 131172 118532 131178 118544
rect 140038 118532 140044 118544
rect 140096 118532 140102 118584
rect 131206 118464 131212 118516
rect 131264 118504 131270 118516
rect 134610 118504 134616 118516
rect 131264 118476 134616 118504
rect 131264 118464 131270 118476
rect 134610 118464 134616 118476
rect 134668 118464 134674 118516
rect 145650 117308 145656 117360
rect 145708 117348 145714 117360
rect 186314 117348 186320 117360
rect 145708 117320 186320 117348
rect 145708 117308 145714 117320
rect 186314 117308 186320 117320
rect 186372 117308 186378 117360
rect 411254 117308 411260 117360
rect 411312 117348 411318 117360
rect 436830 117348 436836 117360
rect 411312 117320 436836 117348
rect 411312 117308 411318 117320
rect 436830 117308 436836 117320
rect 436888 117308 436894 117360
rect 131206 117240 131212 117292
rect 131264 117280 131270 117292
rect 146938 117280 146944 117292
rect 131264 117252 146944 117280
rect 131264 117240 131270 117252
rect 146938 117240 146944 117252
rect 146996 117240 147002 117292
rect 131114 117172 131120 117224
rect 131172 117212 131178 117224
rect 134518 117212 134524 117224
rect 131172 117184 134524 117212
rect 131172 117172 131178 117184
rect 134518 117172 134524 117184
rect 134576 117172 134582 117224
rect 141786 115948 141792 116000
rect 141844 115988 141850 116000
rect 186314 115988 186320 116000
rect 141844 115960 186320 115988
rect 141844 115948 141850 115960
rect 186314 115948 186320 115960
rect 186372 115948 186378 116000
rect 411254 115948 411260 116000
rect 411312 115988 411318 116000
rect 423214 115988 423220 116000
rect 411312 115960 423220 115988
rect 411312 115948 411318 115960
rect 423214 115948 423220 115960
rect 423272 115948 423278 116000
rect 131206 115880 131212 115932
rect 131264 115920 131270 115932
rect 144178 115920 144184 115932
rect 131264 115892 144184 115920
rect 131264 115880 131270 115892
rect 144178 115880 144184 115892
rect 144236 115880 144242 115932
rect 411898 115880 411904 115932
rect 411956 115920 411962 115932
rect 437474 115920 437480 115932
rect 411956 115892 437480 115920
rect 411956 115880 411962 115892
rect 437474 115880 437480 115892
rect 437532 115880 437538 115932
rect 131206 115472 131212 115524
rect 131264 115512 131270 115524
rect 134702 115512 134708 115524
rect 131264 115484 134708 115512
rect 131264 115472 131270 115484
rect 134702 115472 134708 115484
rect 134760 115472 134766 115524
rect 431954 115200 431960 115252
rect 432012 115240 432018 115252
rect 434070 115240 434076 115252
rect 432012 115212 434076 115240
rect 432012 115200 432018 115212
rect 434070 115200 434076 115212
rect 434128 115200 434134 115252
rect 149790 114520 149796 114572
rect 149848 114560 149854 114572
rect 186314 114560 186320 114572
rect 149848 114532 186320 114560
rect 149848 114520 149854 114532
rect 186314 114520 186320 114532
rect 186372 114520 186378 114572
rect 131298 114452 131304 114504
rect 131356 114492 131362 114504
rect 187050 114492 187056 114504
rect 131356 114464 187056 114492
rect 131356 114452 131362 114464
rect 187050 114452 187056 114464
rect 187108 114452 187114 114504
rect 428458 114452 428464 114504
rect 428516 114492 428522 114504
rect 437474 114492 437480 114504
rect 428516 114464 437480 114492
rect 428516 114452 428522 114464
rect 437474 114452 437480 114464
rect 437532 114452 437538 114504
rect 131206 114384 131212 114436
rect 131264 114424 131270 114436
rect 159450 114424 159456 114436
rect 131264 114396 159456 114424
rect 131264 114384 131270 114396
rect 159450 114384 159456 114396
rect 159508 114384 159514 114436
rect 131114 114316 131120 114368
rect 131172 114356 131178 114368
rect 141418 114356 141424 114368
rect 131172 114328 141424 114356
rect 131172 114316 131178 114328
rect 141418 114316 141424 114328
rect 141476 114316 141482 114368
rect 131206 113092 131212 113144
rect 131264 113132 131270 113144
rect 147030 113132 147036 113144
rect 131264 113104 147036 113132
rect 131264 113092 131270 113104
rect 147030 113092 147036 113104
rect 147088 113092 147094 113144
rect 428550 113092 428556 113144
rect 428608 113132 428614 113144
rect 437474 113132 437480 113144
rect 428608 113104 437480 113132
rect 428608 113092 428614 113104
rect 437474 113092 437480 113104
rect 437532 113092 437538 113144
rect 131114 113024 131120 113076
rect 131172 113064 131178 113076
rect 137278 113064 137284 113076
rect 131172 113036 137284 113064
rect 131172 113024 131178 113036
rect 137278 113024 137284 113036
rect 137336 113024 137342 113076
rect 146938 111800 146944 111852
rect 146996 111840 147002 111852
rect 186314 111840 186320 111852
rect 146996 111812 186320 111840
rect 146996 111800 147002 111812
rect 186314 111800 186320 111812
rect 186372 111800 186378 111852
rect 411254 111800 411260 111852
rect 411312 111840 411318 111852
rect 421834 111840 421840 111852
rect 411312 111812 421840 111840
rect 411312 111800 411318 111812
rect 421834 111800 421840 111812
rect 421892 111800 421898 111852
rect 132126 111732 132132 111784
rect 132184 111772 132190 111784
rect 147122 111772 147128 111784
rect 132184 111744 147128 111772
rect 132184 111732 132190 111744
rect 147122 111732 147128 111744
rect 147180 111732 147186 111784
rect 418982 111732 418988 111784
rect 419040 111772 419046 111784
rect 437474 111772 437480 111784
rect 419040 111744 437480 111772
rect 419040 111732 419046 111744
rect 437474 111732 437480 111744
rect 437532 111732 437538 111784
rect 131206 111664 131212 111716
rect 131264 111704 131270 111716
rect 140130 111704 140136 111716
rect 131264 111676 140136 111704
rect 131264 111664 131270 111676
rect 140130 111664 140136 111676
rect 140188 111664 140194 111716
rect 134518 110440 134524 110492
rect 134576 110480 134582 110492
rect 186314 110480 186320 110492
rect 134576 110452 186320 110480
rect 134576 110440 134582 110452
rect 186314 110440 186320 110452
rect 186372 110440 186378 110492
rect 411254 110440 411260 110492
rect 411312 110480 411318 110492
rect 421742 110480 421748 110492
rect 411312 110452 421748 110480
rect 411312 110440 411318 110452
rect 421742 110440 421748 110452
rect 421800 110440 421806 110492
rect 431862 110480 431868 110492
rect 429212 110452 431868 110480
rect 131298 110372 131304 110424
rect 131356 110412 131362 110424
rect 133322 110412 133328 110424
rect 131356 110384 133328 110412
rect 131356 110372 131362 110384
rect 133322 110372 133328 110384
rect 133380 110372 133386 110424
rect 427814 110372 427820 110424
rect 427872 110412 427878 110424
rect 429212 110412 429240 110452
rect 431862 110440 431868 110452
rect 431920 110440 431926 110492
rect 427872 110384 429240 110412
rect 427872 110372 427878 110384
rect 131206 110304 131212 110356
rect 131264 110344 131270 110356
rect 156690 110344 156696 110356
rect 131264 110316 156696 110344
rect 131264 110304 131270 110316
rect 156690 110304 156696 110316
rect 156748 110304 156754 110356
rect 428642 110304 428648 110356
rect 428700 110344 428706 110356
rect 437474 110344 437480 110356
rect 428700 110316 437480 110344
rect 428700 110304 428706 110316
rect 437474 110304 437480 110316
rect 437532 110304 437538 110356
rect 131114 110236 131120 110288
rect 131172 110276 131178 110288
rect 159542 110276 159548 110288
rect 131172 110248 159548 110276
rect 131172 110236 131178 110248
rect 159542 110236 159548 110248
rect 159600 110236 159606 110288
rect 141418 109012 141424 109064
rect 141476 109052 141482 109064
rect 186314 109052 186320 109064
rect 141476 109024 186320 109052
rect 141476 109012 141482 109024
rect 186314 109012 186320 109024
rect 186372 109012 186378 109064
rect 131114 108944 131120 108996
rect 131172 108984 131178 108996
rect 141510 108984 141516 108996
rect 131172 108956 141516 108984
rect 131172 108944 131178 108956
rect 141510 108944 141516 108956
rect 141568 108944 141574 108996
rect 131206 108876 131212 108928
rect 131264 108916 131270 108928
rect 137370 108916 137376 108928
rect 131264 108888 137376 108916
rect 131264 108876 131270 108888
rect 137370 108876 137376 108888
rect 137428 108876 137434 108928
rect 424962 108060 424968 108112
rect 425020 108100 425026 108112
rect 427814 108100 427820 108112
rect 425020 108072 427820 108100
rect 425020 108060 425026 108072
rect 427814 108060 427820 108072
rect 427872 108060 427878 108112
rect 147030 107652 147036 107704
rect 147088 107692 147094 107704
rect 186314 107692 186320 107704
rect 147088 107664 186320 107692
rect 147088 107652 147094 107664
rect 186314 107652 186320 107664
rect 186372 107652 186378 107704
rect 131114 107584 131120 107636
rect 131172 107624 131178 107636
rect 156874 107624 156880 107636
rect 131172 107596 156880 107624
rect 131172 107584 131178 107596
rect 156874 107584 156880 107596
rect 156932 107584 156938 107636
rect 131298 107516 131304 107568
rect 131356 107556 131362 107568
rect 140314 107556 140320 107568
rect 131356 107528 140320 107556
rect 131356 107516 131362 107528
rect 140314 107516 140320 107528
rect 140372 107516 140378 107568
rect 131206 107448 131212 107500
rect 131264 107488 131270 107500
rect 140222 107488 140228 107500
rect 131264 107460 140228 107488
rect 131264 107448 131270 107460
rect 140222 107448 140228 107460
rect 140280 107448 140286 107500
rect 418154 106700 418160 106752
rect 418212 106740 418218 106752
rect 424962 106740 424968 106752
rect 418212 106712 424968 106740
rect 418212 106700 418218 106712
rect 424962 106700 424968 106712
rect 425020 106700 425026 106752
rect 147122 106360 147128 106412
rect 147180 106400 147186 106412
rect 186406 106400 186412 106412
rect 147180 106372 186412 106400
rect 147180 106360 147186 106372
rect 186406 106360 186412 106372
rect 186464 106360 186470 106412
rect 140038 106292 140044 106344
rect 140096 106332 140102 106344
rect 186314 106332 186320 106344
rect 140096 106304 186320 106332
rect 140096 106292 140102 106304
rect 186314 106292 186320 106304
rect 186372 106292 186378 106344
rect 411254 106292 411260 106344
rect 411312 106332 411318 106344
rect 417786 106332 417792 106344
rect 411312 106304 417792 106332
rect 411312 106292 411318 106304
rect 417786 106292 417792 106304
rect 417844 106292 417850 106344
rect 131114 106224 131120 106276
rect 131172 106264 131178 106276
rect 156782 106264 156788 106276
rect 131172 106236 156788 106264
rect 131172 106224 131178 106236
rect 156782 106224 156788 106236
rect 156840 106224 156846 106276
rect 425698 106224 425704 106276
rect 425756 106264 425762 106276
rect 437474 106264 437480 106276
rect 425756 106236 437480 106264
rect 425756 106224 425762 106236
rect 437474 106224 437480 106236
rect 437532 106224 437538 106276
rect 131206 106156 131212 106208
rect 131264 106196 131270 106208
rect 137462 106196 137468 106208
rect 131264 106168 137468 106196
rect 131264 106156 131270 106168
rect 137462 106156 137468 106168
rect 137520 106156 137526 106208
rect 141510 104864 141516 104916
rect 141568 104904 141574 104916
rect 186314 104904 186320 104916
rect 141568 104876 186320 104904
rect 141568 104864 141574 104876
rect 186314 104864 186320 104876
rect 186372 104864 186378 104916
rect 131206 104796 131212 104848
rect 131264 104836 131270 104848
rect 144270 104836 144276 104848
rect 131264 104808 144276 104836
rect 131264 104796 131270 104808
rect 144270 104796 144276 104808
rect 144328 104796 144334 104848
rect 435358 104796 435364 104848
rect 435416 104836 435422 104848
rect 437658 104836 437664 104848
rect 435416 104808 437664 104836
rect 435416 104796 435422 104808
rect 437658 104796 437664 104808
rect 437716 104796 437722 104848
rect 131114 104728 131120 104780
rect 131172 104768 131178 104780
rect 138658 104768 138664 104780
rect 131172 104740 138664 104768
rect 131172 104728 131178 104740
rect 138658 104728 138664 104740
rect 138716 104728 138722 104780
rect 134610 103504 134616 103556
rect 134668 103544 134674 103556
rect 186314 103544 186320 103556
rect 134668 103516 186320 103544
rect 134668 103504 134674 103516
rect 186314 103504 186320 103516
rect 186372 103504 186378 103556
rect 411254 103504 411260 103556
rect 411312 103544 411318 103556
rect 413370 103544 413376 103556
rect 411312 103516 413376 103544
rect 411312 103504 411318 103516
rect 413370 103504 413376 103516
rect 413428 103504 413434 103556
rect 131666 103436 131672 103488
rect 131724 103476 131730 103488
rect 164970 103476 164976 103488
rect 131724 103448 164976 103476
rect 131724 103436 131730 103448
rect 164970 103436 164976 103448
rect 165028 103436 165034 103488
rect 417418 103436 417424 103488
rect 417476 103476 417482 103488
rect 437474 103476 437480 103488
rect 417476 103448 437480 103476
rect 417476 103436 417482 103448
rect 437474 103436 437480 103448
rect 437532 103436 437538 103488
rect 131206 103368 131212 103420
rect 131264 103408 131270 103420
rect 141602 103408 141608 103420
rect 131264 103380 141608 103408
rect 131264 103368 131270 103380
rect 141602 103368 141608 103380
rect 141660 103368 141666 103420
rect 131114 103300 131120 103352
rect 131172 103340 131178 103352
rect 138750 103340 138756 103352
rect 131172 103312 138756 103340
rect 131172 103300 131178 103312
rect 138750 103300 138756 103312
rect 138808 103300 138814 103352
rect 140130 102144 140136 102196
rect 140188 102184 140194 102196
rect 186314 102184 186320 102196
rect 140188 102156 186320 102184
rect 140188 102144 140194 102156
rect 186314 102144 186320 102156
rect 186372 102144 186378 102196
rect 411254 102144 411260 102196
rect 411312 102184 411318 102196
rect 418982 102184 418988 102196
rect 411312 102156 418988 102184
rect 411312 102144 411318 102156
rect 418982 102144 418988 102156
rect 419040 102144 419046 102196
rect 131206 102076 131212 102128
rect 131264 102116 131270 102128
rect 160830 102116 160836 102128
rect 131264 102088 160836 102116
rect 131264 102076 131270 102088
rect 160830 102076 160836 102088
rect 160888 102076 160894 102128
rect 414934 102076 414940 102128
rect 414992 102116 414998 102128
rect 437474 102116 437480 102128
rect 414992 102088 437480 102116
rect 414992 102076 414998 102088
rect 437474 102076 437480 102088
rect 437532 102076 437538 102128
rect 131114 102008 131120 102060
rect 131172 102048 131178 102060
rect 137554 102048 137560 102060
rect 131172 102020 137560 102048
rect 131172 102008 131178 102020
rect 137554 102008 137560 102020
rect 137612 102008 137618 102060
rect 133690 101396 133696 101448
rect 133748 101436 133754 101448
rect 187418 101436 187424 101448
rect 133748 101408 187424 101436
rect 133748 101396 133754 101408
rect 187418 101396 187424 101408
rect 187476 101396 187482 101448
rect 134702 100716 134708 100768
rect 134760 100756 134766 100768
rect 186314 100756 186320 100768
rect 134760 100728 186320 100756
rect 134760 100716 134766 100728
rect 186314 100716 186320 100728
rect 186372 100716 186378 100768
rect 411254 100716 411260 100768
rect 411312 100756 411318 100768
rect 417418 100756 417424 100768
rect 411312 100728 417424 100756
rect 411312 100716 411318 100728
rect 417418 100716 417424 100728
rect 417476 100716 417482 100768
rect 131206 100648 131212 100700
rect 131264 100688 131270 100700
rect 158162 100688 158168 100700
rect 131264 100660 158168 100688
rect 131264 100648 131270 100660
rect 158162 100648 158168 100660
rect 158220 100648 158226 100700
rect 540422 100648 540428 100700
rect 540480 100688 540486 100700
rect 580166 100688 580172 100700
rect 540480 100660 580172 100688
rect 540480 100648 540486 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 131482 99968 131488 100020
rect 131540 100008 131546 100020
rect 159634 100008 159640 100020
rect 131540 99980 159640 100008
rect 131540 99968 131546 99980
rect 159634 99968 159640 99980
rect 159692 99968 159698 100020
rect 144178 99356 144184 99408
rect 144236 99396 144242 99408
rect 186314 99396 186320 99408
rect 144236 99368 186320 99396
rect 144236 99356 144242 99368
rect 186314 99356 186320 99368
rect 186372 99356 186378 99408
rect 415946 99356 415952 99408
rect 416004 99396 416010 99408
rect 417878 99396 417884 99408
rect 416004 99368 417884 99396
rect 416004 99356 416010 99368
rect 417878 99356 417884 99368
rect 417936 99356 417942 99408
rect 131206 99288 131212 99340
rect 131264 99328 131270 99340
rect 162210 99328 162216 99340
rect 131264 99300 162216 99328
rect 131264 99288 131270 99300
rect 162210 99288 162216 99300
rect 162268 99288 162274 99340
rect 432598 99288 432604 99340
rect 432656 99328 432662 99340
rect 437474 99328 437480 99340
rect 432656 99300 437480 99328
rect 432656 99288 432662 99300
rect 437474 99288 437480 99300
rect 437532 99288 437538 99340
rect 131114 99220 131120 99272
rect 131172 99260 131178 99272
rect 158254 99260 158260 99272
rect 131172 99232 158260 99260
rect 131172 99220 131178 99232
rect 158254 99220 158260 99232
rect 158312 99220 158318 99272
rect 141602 98064 141608 98116
rect 141660 98104 141666 98116
rect 186406 98104 186412 98116
rect 141660 98076 186412 98104
rect 141660 98064 141666 98076
rect 186406 98064 186412 98076
rect 186464 98064 186470 98116
rect 131850 97996 131856 98048
rect 131908 98036 131914 98048
rect 186314 98036 186320 98048
rect 131908 98008 186320 98036
rect 131908 97996 131914 98008
rect 186314 97996 186320 98008
rect 186372 97996 186378 98048
rect 411254 97996 411260 98048
rect 411312 98036 411318 98048
rect 414934 98036 414940 98048
rect 411312 98008 414940 98036
rect 411312 97996 411318 98008
rect 414934 97996 414940 98008
rect 414992 97996 414998 98048
rect 131114 97928 131120 97980
rect 131172 97968 131178 97980
rect 160922 97968 160928 97980
rect 131172 97940 160928 97968
rect 131172 97928 131178 97940
rect 160922 97928 160928 97940
rect 160980 97928 160986 97980
rect 431218 97928 431224 97980
rect 431276 97968 431282 97980
rect 437474 97968 437480 97980
rect 431276 97940 437480 97968
rect 431276 97928 431282 97940
rect 437474 97928 437480 97940
rect 437532 97928 437538 97980
rect 131206 97860 131212 97912
rect 131264 97900 131270 97912
rect 155310 97900 155316 97912
rect 131264 97872 155316 97900
rect 131264 97860 131270 97872
rect 155310 97860 155316 97872
rect 155368 97860 155374 97912
rect 140222 96636 140228 96688
rect 140280 96676 140286 96688
rect 186314 96676 186320 96688
rect 140280 96648 186320 96676
rect 140280 96636 140286 96648
rect 186314 96636 186320 96648
rect 186372 96636 186378 96688
rect 131114 96568 131120 96620
rect 131172 96608 131178 96620
rect 158346 96608 158352 96620
rect 131172 96580 158352 96608
rect 131172 96568 131178 96580
rect 158346 96568 158352 96580
rect 158404 96568 158410 96620
rect 429838 96568 429844 96620
rect 429896 96608 429902 96620
rect 437474 96608 437480 96620
rect 429896 96580 437480 96608
rect 429896 96568 429902 96580
rect 437474 96568 437480 96580
rect 437532 96568 437538 96620
rect 131206 96432 131212 96484
rect 131264 96472 131270 96484
rect 134794 96472 134800 96484
rect 131264 96444 134800 96472
rect 131264 96432 131270 96444
rect 134794 96432 134800 96444
rect 134852 96432 134858 96484
rect 414014 96024 414020 96076
rect 414072 96064 414078 96076
rect 415946 96064 415952 96076
rect 414072 96036 415952 96064
rect 414072 96024 414078 96036
rect 415946 96024 415952 96036
rect 416004 96024 416010 96076
rect 132218 95956 132224 96008
rect 132276 95996 132282 96008
rect 133506 95996 133512 96008
rect 132276 95968 133512 95996
rect 132276 95956 132282 95968
rect 133506 95956 133512 95968
rect 133564 95956 133570 96008
rect 140314 95208 140320 95260
rect 140372 95248 140378 95260
rect 186314 95248 186320 95260
rect 140372 95220 186320 95248
rect 140372 95208 140378 95220
rect 186314 95208 186320 95220
rect 186372 95208 186378 95260
rect 131206 95140 131212 95192
rect 131264 95180 131270 95192
rect 156966 95180 156972 95192
rect 131264 95152 156972 95180
rect 131264 95140 131270 95152
rect 156966 95140 156972 95152
rect 157024 95140 157030 95192
rect 428734 95140 428740 95192
rect 428792 95180 428798 95192
rect 437474 95180 437480 95192
rect 428792 95152 437480 95180
rect 428792 95140 428798 95152
rect 437474 95140 437480 95152
rect 437532 95140 437538 95192
rect 131114 95072 131120 95124
rect 131172 95112 131178 95124
rect 133414 95112 133420 95124
rect 131172 95084 133420 95112
rect 131172 95072 131178 95084
rect 133414 95072 133420 95084
rect 133472 95072 133478 95124
rect 131942 93848 131948 93900
rect 132000 93888 132006 93900
rect 186314 93888 186320 93900
rect 132000 93860 186320 93888
rect 132000 93848 132006 93860
rect 186314 93848 186320 93860
rect 186372 93848 186378 93900
rect 131206 93780 131212 93832
rect 131264 93820 131270 93832
rect 136082 93820 136088 93832
rect 131264 93792 136088 93820
rect 131264 93780 131270 93792
rect 136082 93780 136088 93792
rect 136140 93780 136146 93832
rect 425790 93780 425796 93832
rect 425848 93820 425854 93832
rect 437474 93820 437480 93832
rect 425848 93792 437480 93820
rect 425848 93780 425854 93792
rect 437474 93780 437480 93792
rect 437532 93780 437538 93832
rect 131114 93712 131120 93764
rect 131172 93752 131178 93764
rect 133598 93752 133604 93764
rect 131172 93724 133604 93752
rect 131172 93712 131178 93724
rect 133598 93712 133604 93724
rect 133656 93712 133662 93764
rect 133230 92488 133236 92540
rect 133288 92528 133294 92540
rect 186314 92528 186320 92540
rect 133288 92500 186320 92528
rect 133288 92488 133294 92500
rect 186314 92488 186320 92500
rect 186372 92488 186378 92540
rect 411346 92488 411352 92540
rect 411404 92528 411410 92540
rect 435358 92528 435364 92540
rect 411404 92500 435364 92528
rect 411404 92488 411410 92500
rect 435358 92488 435364 92500
rect 435416 92488 435422 92540
rect 131298 92420 131304 92472
rect 131356 92460 131362 92472
rect 166350 92460 166356 92472
rect 131356 92432 166356 92460
rect 131356 92420 131362 92432
rect 166350 92420 166356 92432
rect 166408 92420 166414 92472
rect 411254 92420 411260 92472
rect 411312 92460 411318 92472
rect 421926 92460 421932 92472
rect 411312 92432 421932 92460
rect 411312 92420 411318 92432
rect 421926 92420 421932 92432
rect 421984 92420 421990 92472
rect 131114 92352 131120 92404
rect 131172 92392 131178 92404
rect 141694 92392 141700 92404
rect 131172 92364 141700 92392
rect 131172 92352 131178 92364
rect 141694 92352 141700 92364
rect 141752 92352 141758 92404
rect 131206 92284 131212 92336
rect 131264 92324 131270 92336
rect 138842 92324 138848 92336
rect 131264 92296 138848 92324
rect 131264 92284 131270 92296
rect 138842 92284 138848 92296
rect 138900 92284 138906 92336
rect 181438 91060 181444 91112
rect 181496 91100 181502 91112
rect 186314 91100 186320 91112
rect 181496 91072 186320 91100
rect 181496 91060 181502 91072
rect 186314 91060 186320 91072
rect 186372 91060 186378 91112
rect 414014 91100 414020 91112
rect 412606 91072 414020 91100
rect 131206 90992 131212 91044
rect 131264 91032 131270 91044
rect 155402 91032 155408 91044
rect 131264 91004 155408 91032
rect 131264 90992 131270 91004
rect 155402 90992 155408 91004
rect 155460 90992 155466 91044
rect 410518 90992 410524 91044
rect 410576 91032 410582 91044
rect 412606 91032 412634 91072
rect 414014 91060 414020 91072
rect 414072 91060 414078 91112
rect 410576 91004 412634 91032
rect 410576 90992 410582 91004
rect 424318 90992 424324 91044
rect 424376 91032 424382 91044
rect 437474 91032 437480 91044
rect 424376 91004 437480 91032
rect 424376 90992 424382 91004
rect 437474 90992 437480 91004
rect 437532 90992 437538 91044
rect 131114 90924 131120 90976
rect 131172 90964 131178 90976
rect 151170 90964 151176 90976
rect 131172 90936 151176 90964
rect 131172 90924 131178 90936
rect 151170 90924 151176 90936
rect 151228 90924 151234 90976
rect 415026 90312 415032 90364
rect 415084 90352 415090 90364
rect 438302 90352 438308 90364
rect 415084 90324 438308 90352
rect 415084 90312 415090 90324
rect 438302 90312 438308 90324
rect 438360 90312 438366 90364
rect 133322 89700 133328 89752
rect 133380 89740 133386 89752
rect 186314 89740 186320 89752
rect 133380 89712 186320 89740
rect 133380 89700 133386 89712
rect 186314 89700 186320 89712
rect 186372 89700 186378 89752
rect 131298 89632 131304 89684
rect 131356 89672 131362 89684
rect 155494 89672 155500 89684
rect 131356 89644 155500 89672
rect 131356 89632 131362 89644
rect 155494 89632 155500 89644
rect 155552 89632 155558 89684
rect 411254 89632 411260 89684
rect 411312 89672 411318 89684
rect 413554 89672 413560 89684
rect 411312 89644 413560 89672
rect 411312 89632 411318 89644
rect 413554 89632 413560 89644
rect 413612 89632 413618 89684
rect 424410 89632 424416 89684
rect 424468 89672 424474 89684
rect 437474 89672 437480 89684
rect 424468 89644 437480 89672
rect 424468 89632 424474 89644
rect 437474 89632 437480 89644
rect 437532 89632 437538 89684
rect 132218 89564 132224 89616
rect 132276 89604 132282 89616
rect 144362 89604 144368 89616
rect 132276 89576 144368 89604
rect 132276 89564 132282 89576
rect 144362 89564 144368 89576
rect 144420 89564 144426 89616
rect 131114 88952 131120 89004
rect 131172 88992 131178 89004
rect 144454 88992 144460 89004
rect 131172 88964 144460 88992
rect 131172 88952 131178 88964
rect 144454 88952 144460 88964
rect 144512 88952 144518 89004
rect 411806 88952 411812 89004
rect 411864 88992 411870 89004
rect 412174 88992 412180 89004
rect 411864 88964 412180 88992
rect 411864 88952 411870 88964
rect 412174 88952 412180 88964
rect 412232 88952 412238 89004
rect 138658 88340 138664 88392
rect 138716 88380 138722 88392
rect 186314 88380 186320 88392
rect 138716 88352 186320 88380
rect 138716 88340 138722 88352
rect 186314 88340 186320 88352
rect 186372 88340 186378 88392
rect 131298 88272 131304 88324
rect 131356 88312 131362 88324
rect 152458 88312 152464 88324
rect 131356 88284 152464 88312
rect 131356 88272 131362 88284
rect 152458 88272 152464 88284
rect 152516 88272 152522 88324
rect 411254 88272 411260 88324
rect 411312 88312 411318 88324
rect 439958 88312 439964 88324
rect 411312 88284 439964 88312
rect 411312 88272 411318 88284
rect 439958 88272 439964 88284
rect 440016 88272 440022 88324
rect 131206 88204 131212 88256
rect 131264 88244 131270 88256
rect 151262 88244 151268 88256
rect 131264 88216 151268 88244
rect 131264 88204 131270 88216
rect 151262 88204 151268 88216
rect 151320 88204 151326 88256
rect 423122 88204 423128 88256
rect 423180 88244 423186 88256
rect 437474 88244 437480 88256
rect 423180 88216 437480 88244
rect 423180 88204 423186 88216
rect 437474 88204 437480 88216
rect 437532 88204 437538 88256
rect 132034 86980 132040 87032
rect 132092 87020 132098 87032
rect 186314 87020 186320 87032
rect 132092 86992 186320 87020
rect 132092 86980 132098 86992
rect 186314 86980 186320 86992
rect 186372 86980 186378 87032
rect 131114 86912 131120 86964
rect 131172 86952 131178 86964
rect 187142 86952 187148 86964
rect 131172 86924 187148 86952
rect 131172 86912 131178 86924
rect 187142 86912 187148 86924
rect 187200 86912 187206 86964
rect 411254 86912 411260 86964
rect 411312 86952 411318 86964
rect 439866 86952 439872 86964
rect 411312 86924 439872 86952
rect 411312 86912 411318 86924
rect 439866 86912 439872 86924
rect 439924 86912 439930 86964
rect 131206 86844 131212 86896
rect 131264 86884 131270 86896
rect 148410 86884 148416 86896
rect 131264 86856 148416 86884
rect 131264 86844 131270 86856
rect 148410 86844 148416 86856
rect 148468 86844 148474 86896
rect 425882 86844 425888 86896
rect 425940 86884 425946 86896
rect 437474 86884 437480 86896
rect 425940 86856 437480 86884
rect 425940 86844 425946 86856
rect 437474 86844 437480 86856
rect 437532 86844 437538 86896
rect 133414 85552 133420 85604
rect 133472 85592 133478 85604
rect 186314 85592 186320 85604
rect 133472 85564 186320 85592
rect 133472 85552 133478 85564
rect 186314 85552 186320 85564
rect 186372 85552 186378 85604
rect 540422 85552 540428 85604
rect 540480 85592 540486 85604
rect 580166 85592 580172 85604
rect 540480 85564 580172 85592
rect 540480 85552 540486 85564
rect 580166 85552 580172 85564
rect 580224 85552 580230 85604
rect 132218 85484 132224 85536
rect 132276 85524 132282 85536
rect 152550 85524 152556 85536
rect 132276 85496 152556 85524
rect 132276 85484 132282 85496
rect 152550 85484 152556 85496
rect 152608 85484 152614 85536
rect 423030 85484 423036 85536
rect 423088 85524 423094 85536
rect 437474 85524 437480 85536
rect 423088 85496 437480 85524
rect 423088 85484 423094 85496
rect 437474 85484 437480 85496
rect 437532 85484 437538 85536
rect 131114 85416 131120 85468
rect 131172 85456 131178 85468
rect 148502 85456 148508 85468
rect 131172 85428 148508 85456
rect 131172 85416 131178 85428
rect 148502 85416 148508 85428
rect 148560 85416 148566 85468
rect 132218 84804 132224 84856
rect 132276 84844 132282 84856
rect 142890 84844 142896 84856
rect 132276 84816 142896 84844
rect 132276 84804 132282 84816
rect 142890 84804 142896 84816
rect 142948 84804 142954 84856
rect 131206 84124 131212 84176
rect 131264 84164 131270 84176
rect 152642 84164 152648 84176
rect 131264 84136 152648 84164
rect 131264 84124 131270 84136
rect 152642 84124 152648 84136
rect 152700 84124 152706 84176
rect 131114 84056 131120 84108
rect 131172 84096 131178 84108
rect 148594 84096 148600 84108
rect 131172 84068 148600 84096
rect 131172 84056 131178 84068
rect 148594 84056 148600 84068
rect 148652 84056 148658 84108
rect 142890 82900 142896 82952
rect 142948 82940 142954 82952
rect 186314 82940 186320 82952
rect 142948 82912 186320 82940
rect 142948 82900 142954 82912
rect 186314 82900 186320 82912
rect 186372 82900 186378 82952
rect 135990 82832 135996 82884
rect 136048 82872 136054 82884
rect 186406 82872 186412 82884
rect 136048 82844 186412 82872
rect 136048 82832 136054 82844
rect 186406 82832 186412 82844
rect 186464 82832 186470 82884
rect 411254 82832 411260 82884
rect 411312 82872 411318 82884
rect 438210 82872 438216 82884
rect 411312 82844 438216 82872
rect 411312 82832 411318 82844
rect 438210 82832 438216 82844
rect 438268 82832 438274 82884
rect 131574 82764 131580 82816
rect 131632 82804 131638 82816
rect 187234 82804 187240 82816
rect 131632 82776 187240 82804
rect 131632 82764 131638 82776
rect 187234 82764 187240 82776
rect 187292 82764 187298 82816
rect 417510 82764 417516 82816
rect 417568 82804 417574 82816
rect 437474 82804 437480 82816
rect 417568 82776 437480 82804
rect 417568 82764 417574 82776
rect 437474 82764 437480 82776
rect 437532 82764 437538 82816
rect 131206 82696 131212 82748
rect 131264 82736 131270 82748
rect 152734 82736 152740 82748
rect 131264 82708 152740 82736
rect 131264 82696 131270 82708
rect 152734 82696 152740 82708
rect 152792 82696 152798 82748
rect 132218 81336 132224 81388
rect 132276 81376 132282 81388
rect 148686 81376 148692 81388
rect 132276 81348 148692 81376
rect 132276 81336 132282 81348
rect 148686 81336 148692 81348
rect 148744 81336 148750 81388
rect 422938 81336 422944 81388
rect 422996 81376 423002 81388
rect 437474 81376 437480 81388
rect 422996 81348 437480 81376
rect 422996 81336 423002 81348
rect 437474 81336 437480 81348
rect 437532 81336 437538 81388
rect 131206 81268 131212 81320
rect 131264 81308 131270 81320
rect 142982 81308 142988 81320
rect 131264 81280 142988 81308
rect 131264 81268 131270 81280
rect 142982 81268 142988 81280
rect 143040 81268 143046 81320
rect 411254 80112 411260 80164
rect 411312 80152 411318 80164
rect 413554 80152 413560 80164
rect 411312 80124 413560 80152
rect 411312 80112 411318 80124
rect 413554 80112 413560 80124
rect 413612 80112 413618 80164
rect 136082 80044 136088 80096
rect 136140 80084 136146 80096
rect 186314 80084 186320 80096
rect 136140 80056 186320 80084
rect 136140 80044 136146 80056
rect 186314 80044 186320 80056
rect 186372 80044 186378 80096
rect 131206 79976 131212 80028
rect 131264 80016 131270 80028
rect 151354 80016 151360 80028
rect 131264 79988 151360 80016
rect 131264 79976 131270 79988
rect 151354 79976 151360 79988
rect 151412 79976 151418 80028
rect 417602 79976 417608 80028
rect 417660 80016 417666 80028
rect 437474 80016 437480 80028
rect 417660 79988 437480 80016
rect 417660 79976 417666 79988
rect 437474 79976 437480 79988
rect 437532 79976 437538 80028
rect 131114 79908 131120 79960
rect 131172 79948 131178 79960
rect 147214 79948 147220 79960
rect 131172 79920 147220 79948
rect 131172 79908 131178 79920
rect 147214 79908 147220 79920
rect 147272 79908 147278 79960
rect 131206 79840 131212 79892
rect 131264 79880 131270 79892
rect 143074 79880 143080 79892
rect 131264 79852 143080 79880
rect 131264 79840 131270 79852
rect 143074 79840 143080 79852
rect 143132 79840 143138 79892
rect 138750 78684 138756 78736
rect 138808 78724 138814 78736
rect 186314 78724 186320 78736
rect 138808 78696 186320 78724
rect 138808 78684 138814 78696
rect 186314 78684 186320 78696
rect 186372 78684 186378 78736
rect 131206 78616 131212 78668
rect 131264 78656 131270 78668
rect 151078 78656 151084 78668
rect 131264 78628 151084 78656
rect 131264 78616 131270 78628
rect 151078 78616 151084 78628
rect 151136 78616 151142 78668
rect 421650 78616 421656 78668
rect 421708 78656 421714 78668
rect 437474 78656 437480 78668
rect 421708 78628 437480 78656
rect 421708 78616 421714 78628
rect 437474 78616 437480 78628
rect 437532 78616 437538 78668
rect 131114 78548 131120 78600
rect 131172 78588 131178 78600
rect 145558 78588 145564 78600
rect 131172 78560 145564 78588
rect 131172 78548 131178 78560
rect 145558 78548 145564 78560
rect 145616 78548 145622 78600
rect 411254 78276 411260 78328
rect 411312 78316 411318 78328
rect 413646 78316 413652 78328
rect 411312 78288 413652 78316
rect 411312 78276 411318 78288
rect 413646 78276 413652 78288
rect 413704 78276 413710 78328
rect 131298 77936 131304 77988
rect 131356 77976 131362 77988
rect 187326 77976 187332 77988
rect 131356 77948 187332 77976
rect 131356 77936 131362 77948
rect 187326 77936 187332 77948
rect 187384 77936 187390 77988
rect 131206 77188 131212 77240
rect 131264 77228 131270 77240
rect 149698 77228 149704 77240
rect 131264 77200 149704 77228
rect 131264 77188 131270 77200
rect 149698 77188 149704 77200
rect 149756 77188 149762 77240
rect 411254 77188 411260 77240
rect 411312 77228 411318 77240
rect 438118 77228 438124 77240
rect 411312 77200 438124 77228
rect 411312 77188 411318 77200
rect 438118 77188 438124 77200
rect 438176 77188 438182 77240
rect 131114 77120 131120 77172
rect 131172 77160 131178 77172
rect 145742 77160 145748 77172
rect 131172 77132 145748 77160
rect 131172 77120 131178 77132
rect 145742 77120 145748 77132
rect 145800 77120 145806 77172
rect 138842 75964 138848 76016
rect 138900 76004 138906 76016
rect 186314 76004 186320 76016
rect 138900 75976 186320 76004
rect 138900 75964 138906 75976
rect 186314 75964 186320 75976
rect 186372 75964 186378 76016
rect 134794 75896 134800 75948
rect 134852 75936 134858 75948
rect 186406 75936 186412 75948
rect 134852 75908 186412 75936
rect 134852 75896 134858 75908
rect 186406 75896 186412 75908
rect 186464 75896 186470 75948
rect 131206 75828 131212 75880
rect 131264 75868 131270 75880
rect 142798 75868 142804 75880
rect 131264 75840 142804 75868
rect 131264 75828 131270 75840
rect 142798 75828 142804 75840
rect 142856 75828 142862 75880
rect 419166 75828 419172 75880
rect 419224 75868 419230 75880
rect 437474 75868 437480 75880
rect 419224 75840 437480 75868
rect 419224 75828 419230 75840
rect 437474 75828 437480 75840
rect 437532 75828 437538 75880
rect 131114 75760 131120 75812
rect 131172 75800 131178 75812
rect 135898 75800 135904 75812
rect 131172 75772 135904 75800
rect 131172 75760 131178 75772
rect 135898 75760 135904 75772
rect 135956 75760 135962 75812
rect 159358 75216 159364 75268
rect 159416 75256 159422 75268
rect 187510 75256 187516 75268
rect 159416 75228 187516 75256
rect 159416 75216 159422 75228
rect 187510 75216 187516 75228
rect 187568 75216 187574 75268
rect 132494 75148 132500 75200
rect 132552 75188 132558 75200
rect 186958 75188 186964 75200
rect 132552 75160 186964 75188
rect 132552 75148 132558 75160
rect 186958 75148 186964 75160
rect 187016 75148 187022 75200
rect 131206 74468 131212 74520
rect 131264 74508 131270 74520
rect 145650 74508 145656 74520
rect 131264 74480 145656 74508
rect 131264 74468 131270 74480
rect 145650 74468 145656 74480
rect 145708 74468 145714 74520
rect 411254 74468 411260 74520
rect 411312 74508 411318 74520
rect 435542 74508 435548 74520
rect 411312 74480 435548 74508
rect 411312 74468 411318 74480
rect 435542 74468 435548 74480
rect 435600 74468 435606 74520
rect 131114 74400 131120 74452
rect 131172 74440 131178 74452
rect 141786 74440 141792 74452
rect 131172 74412 141792 74440
rect 131172 74400 131178 74412
rect 141786 74400 141792 74412
rect 141844 74400 141850 74452
rect 421558 74400 421564 74452
rect 421616 74440 421622 74452
rect 437474 74440 437480 74452
rect 421616 74412 437480 74440
rect 421616 74400 421622 74412
rect 437474 74400 437480 74412
rect 437532 74400 437538 74452
rect 132310 73176 132316 73228
rect 132368 73216 132374 73228
rect 186314 73216 186320 73228
rect 132368 73188 186320 73216
rect 132368 73176 132374 73188
rect 186314 73176 186320 73188
rect 186372 73176 186378 73228
rect 131114 73108 131120 73160
rect 131172 73148 131178 73160
rect 133690 73148 133696 73160
rect 131172 73120 133696 73148
rect 131172 73108 131178 73120
rect 133690 73108 133696 73120
rect 133748 73108 133754 73160
rect 429930 73108 429936 73160
rect 429988 73148 429994 73160
rect 437474 73148 437480 73160
rect 429988 73120 437480 73148
rect 429988 73108 429994 73120
rect 437474 73108 437480 73120
rect 437532 73108 437538 73160
rect 131206 72972 131212 73024
rect 131264 73012 131270 73024
rect 149790 73012 149796 73024
rect 131264 72984 149796 73012
rect 131264 72972 131270 72984
rect 149790 72972 149796 72984
rect 149848 72972 149854 73024
rect 411254 72768 411260 72820
rect 411312 72808 411318 72820
rect 413462 72808 413468 72820
rect 411312 72780 413468 72808
rect 411312 72768 411318 72780
rect 413462 72768 413468 72780
rect 413520 72768 413526 72820
rect 181530 71748 181536 71800
rect 181588 71788 181594 71800
rect 186314 71788 186320 71800
rect 181588 71760 186320 71788
rect 181588 71748 181594 71760
rect 186314 71748 186320 71760
rect 186372 71748 186378 71800
rect 131206 71680 131212 71732
rect 131264 71720 131270 71732
rect 146938 71720 146944 71732
rect 131264 71692 146944 71720
rect 131264 71680 131270 71692
rect 146938 71680 146944 71692
rect 146996 71680 147002 71732
rect 417694 71680 417700 71732
rect 417752 71720 417758 71732
rect 437474 71720 437480 71732
rect 417752 71692 437480 71720
rect 417752 71680 417758 71692
rect 437474 71680 437480 71692
rect 437532 71680 437538 71732
rect 131114 71612 131120 71664
rect 131172 71652 131178 71664
rect 134518 71652 134524 71664
rect 131172 71624 134524 71652
rect 131172 71612 131178 71624
rect 134518 71612 134524 71624
rect 134576 71612 134582 71664
rect 133506 70388 133512 70440
rect 133564 70428 133570 70440
rect 186314 70428 186320 70440
rect 133564 70400 186320 70428
rect 133564 70388 133570 70400
rect 186314 70388 186320 70400
rect 186372 70388 186378 70440
rect 131114 70320 131120 70372
rect 131172 70360 131178 70372
rect 147030 70360 147036 70372
rect 131172 70332 147036 70360
rect 131172 70320 131178 70332
rect 147030 70320 147036 70332
rect 147088 70320 147094 70372
rect 426066 70320 426072 70372
rect 426124 70360 426130 70372
rect 437474 70360 437480 70372
rect 426124 70332 437480 70360
rect 426124 70320 426130 70332
rect 437474 70320 437480 70332
rect 437532 70320 437538 70372
rect 131206 70252 131212 70304
rect 131264 70292 131270 70304
rect 141418 70292 141424 70304
rect 131264 70264 141424 70292
rect 131264 70252 131270 70264
rect 141418 70252 141424 70264
rect 141476 70252 141482 70304
rect 146938 69096 146944 69148
rect 146996 69136 147002 69148
rect 186406 69136 186412 69148
rect 146996 69108 186412 69136
rect 146996 69096 147002 69108
rect 186406 69096 186412 69108
rect 186464 69096 186470 69148
rect 134518 69028 134524 69080
rect 134576 69068 134582 69080
rect 186314 69068 186320 69080
rect 134576 69040 186320 69068
rect 134576 69028 134582 69040
rect 186314 69028 186320 69040
rect 186372 69028 186378 69080
rect 131114 68960 131120 69012
rect 131172 69000 131178 69012
rect 147122 69000 147128 69012
rect 131172 68972 147128 69000
rect 131172 68960 131178 68972
rect 147122 68960 147128 68972
rect 147180 68960 147186 69012
rect 131298 68892 131304 68944
rect 131356 68932 131362 68944
rect 141510 68932 141516 68944
rect 131356 68904 141516 68932
rect 131356 68892 131362 68904
rect 141510 68892 141516 68904
rect 141568 68892 141574 68944
rect 131206 68824 131212 68876
rect 131264 68864 131270 68876
rect 140038 68864 140044 68876
rect 131264 68836 140044 68864
rect 131264 68824 131270 68836
rect 140038 68824 140044 68836
rect 140096 68824 140102 68876
rect 181622 67600 181628 67652
rect 181680 67640 181686 67652
rect 186314 67640 186320 67652
rect 181680 67612 186320 67640
rect 181680 67600 181686 67612
rect 186314 67600 186320 67612
rect 186372 67600 186378 67652
rect 411346 67600 411352 67652
rect 411404 67640 411410 67652
rect 439866 67640 439872 67652
rect 411404 67612 439872 67640
rect 411404 67600 411410 67612
rect 439866 67600 439872 67612
rect 439924 67600 439930 67652
rect 131114 67532 131120 67584
rect 131172 67572 131178 67584
rect 140130 67572 140136 67584
rect 131172 67544 140136 67572
rect 131172 67532 131178 67544
rect 140130 67532 140136 67544
rect 140188 67532 140194 67584
rect 411254 67532 411260 67584
rect 411312 67572 411318 67584
rect 439774 67572 439780 67584
rect 411312 67544 439780 67572
rect 411312 67532 411318 67544
rect 439774 67532 439780 67544
rect 439832 67532 439838 67584
rect 425974 67464 425980 67516
rect 426032 67504 426038 67516
rect 437474 67504 437480 67516
rect 426032 67476 437480 67504
rect 426032 67464 426038 67476
rect 437474 67464 437480 67476
rect 437532 67464 437538 67516
rect 131206 67328 131212 67380
rect 131264 67368 131270 67380
rect 134610 67368 134616 67380
rect 131264 67340 134616 67368
rect 131264 67328 131270 67340
rect 134610 67328 134616 67340
rect 134668 67328 134674 67380
rect 144270 66240 144276 66292
rect 144328 66280 144334 66292
rect 186314 66280 186320 66292
rect 144328 66252 186320 66280
rect 144328 66240 144334 66252
rect 186314 66240 186320 66252
rect 186372 66240 186378 66292
rect 131114 66172 131120 66224
rect 131172 66212 131178 66224
rect 144178 66212 144184 66224
rect 131172 66184 144184 66212
rect 131172 66172 131178 66184
rect 144178 66172 144184 66184
rect 144236 66172 144242 66224
rect 431310 66172 431316 66224
rect 431368 66212 431374 66224
rect 437474 66212 437480 66224
rect 431368 66184 437480 66212
rect 431368 66172 431374 66184
rect 437474 66172 437480 66184
rect 437532 66172 437538 66224
rect 131206 66104 131212 66156
rect 131264 66144 131270 66156
rect 134702 66144 134708 66156
rect 131264 66116 134708 66144
rect 131264 66104 131270 66116
rect 134702 66104 134708 66116
rect 134760 66104 134766 66156
rect 411254 65016 411260 65068
rect 411312 65056 411318 65068
rect 413462 65056 413468 65068
rect 411312 65028 413468 65056
rect 411312 65016 411318 65028
rect 413462 65016 413468 65028
rect 413520 65016 413526 65068
rect 134610 64880 134616 64932
rect 134668 64920 134674 64932
rect 186314 64920 186320 64932
rect 134668 64892 186320 64920
rect 134668 64880 134674 64892
rect 186314 64880 186320 64892
rect 186372 64880 186378 64932
rect 131206 64812 131212 64864
rect 131264 64852 131270 64864
rect 141602 64852 141608 64864
rect 131264 64824 141608 64852
rect 131264 64812 131270 64824
rect 141602 64812 141608 64824
rect 141660 64812 141666 64864
rect 424502 64812 424508 64864
rect 424560 64852 424566 64864
rect 437474 64852 437480 64864
rect 424560 64824 437480 64852
rect 424560 64812 424566 64824
rect 437474 64812 437480 64824
rect 437532 64812 437538 64864
rect 131114 64744 131120 64796
rect 131172 64784 131178 64796
rect 140222 64784 140228 64796
rect 131172 64756 140228 64784
rect 131172 64744 131178 64756
rect 140222 64744 140228 64756
rect 140280 64744 140286 64796
rect 181806 63520 181812 63572
rect 181864 63560 181870 63572
rect 186314 63560 186320 63572
rect 181864 63532 186320 63560
rect 181864 63520 181870 63532
rect 186314 63520 186320 63532
rect 186372 63520 186378 63572
rect 132218 63452 132224 63504
rect 132276 63492 132282 63504
rect 140314 63492 140320 63504
rect 132276 63464 140320 63492
rect 132276 63452 132282 63464
rect 140314 63452 140320 63464
rect 140372 63452 140378 63504
rect 411254 63452 411260 63504
rect 411312 63492 411318 63504
rect 420270 63492 420276 63504
rect 411312 63464 420276 63492
rect 411312 63452 411318 63464
rect 420270 63452 420276 63464
rect 420328 63452 420334 63504
rect 142798 62092 142804 62144
rect 142856 62132 142862 62144
rect 186314 62132 186320 62144
rect 142856 62104 186320 62132
rect 142856 62092 142862 62104
rect 186314 62092 186320 62104
rect 186372 62092 186378 62144
rect 131206 62024 131212 62076
rect 131264 62064 131270 62076
rect 133230 62064 133236 62076
rect 131264 62036 133236 62064
rect 131264 62024 131270 62036
rect 133230 62024 133236 62036
rect 133288 62024 133294 62076
rect 424594 62024 424600 62076
rect 424652 62064 424658 62076
rect 437474 62064 437480 62076
rect 424652 62036 437480 62064
rect 424652 62024 424658 62036
rect 437474 62024 437480 62036
rect 437532 62024 437538 62076
rect 132126 61956 132132 62008
rect 132184 61996 132190 62008
rect 159358 61996 159364 62008
rect 132184 61968 159364 61996
rect 132184 61956 132190 61968
rect 159358 61956 159364 61968
rect 159416 61956 159422 62008
rect 131114 61888 131120 61940
rect 131172 61928 131178 61940
rect 181438 61928 181444 61940
rect 131172 61900 181444 61928
rect 131172 61888 131178 61900
rect 181438 61888 181444 61900
rect 181496 61888 181502 61940
rect 181714 60800 181720 60852
rect 181772 60840 181778 60852
rect 186314 60840 186320 60852
rect 181772 60812 186320 60840
rect 181772 60800 181778 60812
rect 186314 60800 186320 60812
rect 186372 60800 186378 60852
rect 134702 60732 134708 60784
rect 134760 60772 134766 60784
rect 186406 60772 186412 60784
rect 134760 60744 186412 60772
rect 134760 60732 134766 60744
rect 186406 60732 186412 60744
rect 186464 60732 186470 60784
rect 411254 60732 411260 60784
rect 411312 60772 411318 60784
rect 439774 60772 439780 60784
rect 411312 60744 439780 60772
rect 411312 60732 411318 60744
rect 439774 60732 439780 60744
rect 439832 60732 439838 60784
rect 131666 60664 131672 60716
rect 131724 60704 131730 60716
rect 138658 60704 138664 60716
rect 131724 60676 138664 60704
rect 131724 60664 131730 60676
rect 138658 60664 138664 60676
rect 138716 60664 138722 60716
rect 411346 60664 411352 60716
rect 411404 60704 411410 60716
rect 420178 60704 420184 60716
rect 411404 60676 420184 60704
rect 411404 60664 411410 60676
rect 420178 60664 420184 60676
rect 420236 60664 420242 60716
rect 540330 60664 540336 60716
rect 540388 60704 540394 60716
rect 580166 60704 580172 60716
rect 540388 60676 580172 60704
rect 540388 60664 540394 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 132218 60596 132224 60648
rect 132276 60636 132282 60648
rect 133322 60636 133328 60648
rect 132276 60608 133328 60636
rect 132276 60596 132282 60608
rect 133322 60596 133328 60608
rect 133380 60596 133386 60648
rect 141418 59372 141424 59424
rect 141476 59412 141482 59424
rect 186314 59412 186320 59424
rect 141476 59384 186320 59412
rect 141476 59372 141482 59384
rect 186314 59372 186320 59384
rect 186372 59372 186378 59424
rect 131298 59304 131304 59356
rect 131356 59344 131362 59356
rect 133414 59344 133420 59356
rect 131356 59316 133420 59344
rect 131356 59304 131362 59316
rect 133414 59304 133420 59316
rect 133472 59304 133478 59356
rect 432690 59304 432696 59356
rect 432748 59344 432754 59356
rect 437474 59344 437480 59356
rect 432748 59316 437480 59344
rect 432748 59304 432754 59316
rect 437474 59304 437480 59316
rect 437532 59304 437538 59356
rect 133230 57944 133236 57996
rect 133288 57984 133294 57996
rect 186314 57984 186320 57996
rect 133288 57956 186320 57984
rect 133288 57944 133294 57956
rect 186314 57944 186320 57956
rect 186372 57944 186378 57996
rect 131206 57876 131212 57928
rect 131264 57916 131270 57928
rect 187050 57916 187056 57928
rect 131264 57888 187056 57916
rect 131264 57876 131270 57888
rect 187050 57876 187056 57888
rect 187108 57876 187114 57928
rect 416038 57876 416044 57928
rect 416096 57916 416102 57928
rect 437474 57916 437480 57928
rect 416096 57888 437480 57916
rect 416096 57876 416102 57888
rect 437474 57876 437480 57888
rect 437532 57876 437538 57928
rect 131114 57808 131120 57860
rect 131172 57848 131178 57860
rect 142890 57848 142896 57860
rect 131172 57820 142896 57848
rect 131172 57808 131178 57820
rect 142890 57808 142896 57820
rect 142948 57808 142954 57860
rect 411254 57808 411260 57860
rect 411312 57848 411318 57860
rect 419074 57848 419080 57860
rect 411312 57820 419080 57848
rect 411312 57808 411318 57820
rect 419074 57808 419080 57820
rect 419132 57808 419138 57860
rect 131206 57740 131212 57792
rect 131264 57780 131270 57792
rect 135990 57780 135996 57792
rect 131264 57752 135996 57780
rect 131264 57740 131270 57752
rect 135990 57740 135996 57752
rect 136048 57740 136054 57792
rect 132218 56516 132224 56568
rect 132276 56556 132282 56568
rect 187142 56556 187148 56568
rect 132276 56528 187148 56556
rect 132276 56516 132282 56528
rect 187142 56516 187148 56528
rect 187200 56516 187206 56568
rect 435450 56516 435456 56568
rect 435508 56556 435514 56568
rect 437750 56556 437756 56568
rect 435508 56528 437756 56556
rect 435508 56516 435514 56528
rect 437750 56516 437756 56528
rect 437808 56516 437814 56568
rect 131206 56448 131212 56500
rect 131264 56488 131270 56500
rect 136082 56488 136088 56500
rect 131264 56460 136088 56488
rect 131264 56448 131270 56460
rect 136082 56448 136088 56460
rect 136140 56448 136146 56500
rect 132494 55836 132500 55888
rect 132552 55876 132558 55888
rect 187418 55876 187424 55888
rect 132552 55848 187424 55876
rect 132552 55836 132558 55848
rect 187418 55836 187424 55848
rect 187476 55836 187482 55888
rect 140038 55224 140044 55276
rect 140096 55264 140102 55276
rect 186314 55264 186320 55276
rect 140096 55236 186320 55264
rect 140096 55224 140102 55236
rect 186314 55224 186320 55236
rect 186372 55224 186378 55276
rect 411254 55224 411260 55276
rect 411312 55264 411318 55276
rect 439958 55264 439964 55276
rect 411312 55236 439964 55264
rect 411312 55224 411318 55236
rect 439958 55224 439964 55236
rect 440016 55224 440022 55276
rect 131206 55156 131212 55208
rect 131264 55196 131270 55208
rect 138750 55196 138756 55208
rect 131264 55168 138756 55196
rect 131264 55156 131270 55168
rect 138750 55156 138756 55168
rect 138808 55156 138814 55208
rect 416130 55156 416136 55208
rect 416188 55196 416194 55208
rect 437474 55196 437480 55208
rect 416188 55168 437480 55196
rect 416188 55156 416194 55168
rect 437474 55156 437480 55168
rect 437532 55156 437538 55208
rect 131298 55088 131304 55140
rect 131356 55128 131362 55140
rect 134794 55128 134800 55140
rect 131356 55100 134800 55128
rect 131356 55088 131362 55100
rect 134794 55088 134800 55100
rect 134852 55088 134858 55140
rect 133322 53796 133328 53848
rect 133380 53836 133386 53848
rect 186314 53836 186320 53848
rect 133380 53808 186320 53836
rect 133380 53796 133386 53808
rect 186314 53796 186320 53808
rect 186372 53796 186378 53848
rect 131114 53728 131120 53780
rect 131172 53768 131178 53780
rect 187234 53768 187240 53780
rect 131172 53740 187240 53768
rect 131172 53728 131178 53740
rect 187234 53728 187240 53740
rect 187292 53728 187298 53780
rect 424686 53728 424692 53780
rect 424744 53768 424750 53780
rect 437474 53768 437480 53780
rect 424744 53740 437480 53768
rect 424744 53728 424750 53740
rect 437474 53728 437480 53740
rect 437532 53728 437538 53780
rect 131206 53660 131212 53712
rect 131264 53700 131270 53712
rect 138842 53700 138848 53712
rect 131264 53672 138848 53700
rect 131264 53660 131270 53672
rect 138842 53660 138848 53672
rect 138900 53660 138906 53712
rect 131850 52436 131856 52488
rect 131908 52476 131914 52488
rect 186314 52476 186320 52488
rect 131908 52448 186320 52476
rect 131908 52436 131914 52448
rect 186314 52436 186320 52448
rect 186372 52436 186378 52488
rect 131206 52368 131212 52420
rect 131264 52408 131270 52420
rect 181530 52408 181536 52420
rect 131264 52380 181536 52408
rect 131264 52368 131270 52380
rect 181530 52368 181536 52380
rect 181588 52368 181594 52420
rect 133414 51076 133420 51128
rect 133472 51116 133478 51128
rect 186314 51116 186320 51128
rect 133472 51088 186320 51116
rect 133472 51076 133478 51088
rect 186314 51076 186320 51088
rect 186372 51076 186378 51128
rect 131114 51008 131120 51060
rect 131172 51048 131178 51060
rect 146938 51048 146944 51060
rect 131172 51020 146944 51048
rect 131172 51008 131178 51020
rect 146938 51008 146944 51020
rect 146996 51008 147002 51060
rect 131206 50940 131212 50992
rect 131264 50980 131270 50992
rect 133506 50980 133512 50992
rect 131264 50952 133512 50980
rect 131264 50940 131270 50952
rect 133506 50940 133512 50952
rect 133564 50940 133570 50992
rect 411254 50940 411260 50992
rect 411312 50980 411318 50992
rect 414750 50980 414756 50992
rect 411312 50952 414756 50980
rect 411312 50940 411318 50952
rect 414750 50940 414756 50952
rect 414808 50940 414814 50992
rect 131298 50872 131304 50924
rect 131356 50912 131362 50924
rect 134518 50912 134524 50924
rect 131356 50884 134524 50912
rect 131356 50872 131362 50884
rect 134518 50872 134524 50884
rect 134576 50872 134582 50924
rect 131206 49648 131212 49700
rect 131264 49688 131270 49700
rect 181622 49688 181628 49700
rect 131264 49660 181628 49688
rect 131264 49648 131270 49660
rect 181622 49648 181628 49660
rect 181680 49648 181686 49700
rect 423214 49648 423220 49700
rect 423272 49688 423278 49700
rect 437474 49688 437480 49700
rect 423272 49660 437480 49688
rect 423272 49648 423278 49660
rect 437474 49648 437480 49660
rect 437532 49648 437538 49700
rect 131114 49580 131120 49632
rect 131172 49620 131178 49632
rect 144270 49620 144276 49632
rect 131172 49592 144276 49620
rect 131172 49580 131178 49592
rect 144270 49580 144276 49592
rect 144328 49580 144334 49632
rect 132034 48288 132040 48340
rect 132092 48328 132098 48340
rect 186314 48328 186320 48340
rect 132092 48300 186320 48328
rect 132092 48288 132098 48300
rect 186314 48288 186320 48300
rect 186372 48288 186378 48340
rect 131206 48220 131212 48272
rect 131264 48260 131270 48272
rect 181806 48260 181812 48272
rect 131264 48232 181812 48260
rect 131264 48220 131270 48232
rect 181806 48220 181812 48232
rect 181864 48220 181870 48272
rect 411990 48220 411996 48272
rect 412048 48260 412054 48272
rect 437474 48260 437480 48272
rect 412048 48232 437480 48260
rect 412048 48220 412054 48232
rect 437474 48220 437480 48232
rect 437532 48220 437538 48272
rect 131942 48016 131948 48068
rect 132000 48056 132006 48068
rect 134610 48056 134616 48068
rect 132000 48028 134616 48056
rect 132000 48016 132006 48028
rect 134610 48016 134616 48028
rect 134668 48016 134674 48068
rect 411254 48016 411260 48068
rect 411312 48056 411318 48068
rect 414842 48056 414848 48068
rect 411312 48028 414848 48056
rect 411312 48016 411318 48028
rect 414842 48016 414848 48028
rect 414900 48016 414906 48068
rect 132494 46928 132500 46980
rect 132552 46968 132558 46980
rect 186314 46968 186320 46980
rect 132552 46940 186320 46968
rect 132552 46928 132558 46940
rect 186314 46928 186320 46940
rect 186372 46928 186378 46980
rect 131206 46860 131212 46912
rect 131264 46900 131270 46912
rect 142798 46900 142804 46912
rect 131264 46872 142804 46900
rect 131264 46860 131270 46872
rect 142798 46860 142804 46872
rect 142856 46860 142862 46912
rect 421834 46860 421840 46912
rect 421892 46900 421898 46912
rect 437474 46900 437480 46912
rect 421892 46872 437480 46900
rect 421892 46860 421898 46872
rect 437474 46860 437480 46872
rect 437532 46860 437538 46912
rect 131114 46792 131120 46844
rect 131172 46832 131178 46844
rect 134702 46832 134708 46844
rect 131172 46804 134708 46832
rect 131172 46792 131178 46804
rect 134702 46792 134708 46804
rect 134760 46792 134766 46844
rect 411254 45568 411260 45620
rect 411312 45608 411318 45620
rect 440050 45608 440056 45620
rect 411312 45580 440056 45608
rect 411312 45568 411318 45580
rect 440050 45568 440056 45580
rect 440108 45568 440114 45620
rect 540330 45568 540336 45620
rect 540388 45608 540394 45620
rect 580166 45608 580172 45620
rect 540388 45580 580172 45608
rect 540388 45568 540394 45580
rect 580166 45568 580172 45580
rect 580224 45568 580230 45620
rect 131298 45500 131304 45552
rect 131356 45540 131362 45552
rect 133230 45540 133236 45552
rect 131356 45512 133236 45540
rect 131356 45500 131362 45512
rect 133230 45500 133236 45512
rect 133288 45500 133294 45552
rect 421742 45500 421748 45552
rect 421800 45540 421806 45552
rect 437474 45540 437480 45552
rect 421800 45512 437480 45540
rect 421800 45500 421806 45512
rect 437474 45500 437480 45512
rect 437532 45500 437538 45552
rect 131114 45432 131120 45484
rect 131172 45472 131178 45484
rect 141418 45472 141424 45484
rect 131172 45444 141424 45472
rect 131172 45432 131178 45444
rect 141418 45432 141424 45444
rect 141476 45432 141482 45484
rect 131206 45364 131212 45416
rect 131264 45404 131270 45416
rect 181714 45404 181720 45416
rect 131264 45376 181720 45404
rect 131264 45364 131270 45376
rect 181714 45364 181720 45376
rect 181772 45364 181778 45416
rect 182082 44140 182088 44192
rect 182140 44180 182146 44192
rect 186314 44180 186320 44192
rect 182140 44152 186320 44180
rect 182140 44140 182146 44152
rect 186314 44140 186320 44152
rect 186372 44140 186378 44192
rect 131206 44072 131212 44124
rect 131264 44112 131270 44124
rect 186958 44112 186964 44124
rect 131264 44084 186964 44112
rect 131264 44072 131270 44084
rect 186958 44072 186964 44084
rect 187016 44072 187022 44124
rect 131114 44004 131120 44056
rect 131172 44044 131178 44056
rect 140038 44044 140044 44056
rect 131172 44016 140044 44044
rect 131172 44004 131178 44016
rect 140038 44004 140044 44016
rect 140096 44004 140102 44056
rect 131298 42780 131304 42832
rect 131356 42820 131362 42832
rect 186314 42820 186320 42832
rect 131356 42792 186320 42820
rect 131356 42780 131362 42792
rect 186314 42780 186320 42792
rect 186372 42780 186378 42832
rect 131114 42712 131120 42764
rect 131172 42752 131178 42764
rect 187050 42752 187056 42764
rect 131172 42724 187056 42752
rect 131172 42712 131178 42724
rect 187050 42712 187056 42724
rect 187108 42712 187114 42764
rect 411898 42712 411904 42764
rect 411956 42752 411962 42764
rect 437474 42752 437480 42764
rect 411956 42724 437480 42752
rect 411956 42712 411962 42724
rect 437474 42712 437480 42724
rect 437532 42712 437538 42764
rect 131206 42644 131212 42696
rect 131264 42684 131270 42696
rect 133322 42684 133328 42696
rect 131264 42656 133328 42684
rect 131264 42644 131270 42656
rect 133322 42644 133328 42656
rect 133380 42644 133386 42696
rect 411254 42508 411260 42560
rect 411312 42548 411318 42560
rect 414658 42548 414664 42560
rect 411312 42520 414664 42548
rect 411312 42508 411318 42520
rect 414658 42508 414664 42520
rect 414716 42508 414722 42560
rect 131114 41352 131120 41404
rect 131172 41392 131178 41404
rect 187142 41392 187148 41404
rect 131172 41364 187148 41392
rect 131172 41352 131178 41364
rect 187142 41352 187148 41364
rect 187200 41352 187206 41404
rect 411254 41352 411260 41404
rect 411312 41392 411318 41404
rect 439682 41392 439688 41404
rect 411312 41364 439688 41392
rect 411312 41352 411318 41364
rect 439682 41352 439688 41364
rect 439740 41352 439746 41404
rect 131206 41284 131212 41336
rect 131264 41324 131270 41336
rect 133414 41324 133420 41336
rect 131264 41296 133420 41324
rect 131264 41284 131270 41296
rect 133414 41284 133420 41296
rect 133472 41284 133478 41336
rect 417786 41284 417792 41336
rect 417844 41324 417850 41336
rect 437474 41324 437480 41336
rect 417844 41296 437480 41324
rect 417844 41284 417850 41296
rect 437474 41284 437480 41296
rect 437532 41284 437538 41336
rect 413370 39992 413376 40044
rect 413428 40032 413434 40044
rect 437474 40032 437480 40044
rect 413428 40004 437480 40032
rect 413428 39992 413434 40004
rect 437474 39992 437480 40004
rect 437532 39992 437538 40044
rect 131482 39312 131488 39364
rect 131540 39352 131546 39364
rect 182082 39352 182088 39364
rect 131540 39324 182088 39352
rect 131540 39312 131546 39324
rect 182082 39312 182088 39324
rect 182140 39312 182146 39364
rect 131850 38632 131856 38684
rect 131908 38672 131914 38684
rect 186314 38672 186320 38684
rect 131908 38644 186320 38672
rect 131908 38632 131914 38644
rect 186314 38632 186320 38644
rect 186372 38632 186378 38684
rect 131206 38564 131212 38616
rect 131264 38604 131270 38616
rect 187418 38604 187424 38616
rect 131264 38576 187424 38604
rect 131264 38564 131270 38576
rect 187418 38564 187424 38576
rect 187476 38564 187482 38616
rect 411254 38564 411260 38616
rect 411312 38604 411318 38616
rect 413278 38604 413284 38616
rect 411312 38576 413284 38604
rect 411312 38564 411318 38576
rect 413278 38564 413284 38576
rect 413336 38564 413342 38616
rect 418982 38564 418988 38616
rect 419040 38604 419046 38616
rect 437474 38604 437480 38616
rect 419040 38576 437480 38604
rect 419040 38564 419046 38576
rect 437474 38564 437480 38576
rect 437532 38564 437538 38616
rect 131114 38496 131120 38548
rect 131172 38536 131178 38548
rect 187234 38536 187240 38548
rect 131172 38508 187240 38536
rect 131172 38496 131178 38508
rect 187234 38496 187240 38508
rect 187292 38496 187298 38548
rect 132126 37272 132132 37324
rect 132184 37312 132190 37324
rect 186314 37312 186320 37324
rect 132184 37284 186320 37312
rect 132184 37272 132190 37284
rect 186314 37272 186320 37284
rect 186372 37272 186378 37324
rect 131206 37204 131212 37256
rect 131264 37244 131270 37256
rect 186406 37244 186412 37256
rect 131264 37216 186412 37244
rect 131264 37204 131270 37216
rect 186406 37204 186412 37216
rect 186464 37204 186470 37256
rect 411254 37204 411260 37256
rect 411312 37244 411318 37256
rect 439590 37244 439596 37256
rect 411312 37216 439596 37244
rect 411312 37204 411318 37216
rect 439590 37204 439596 37216
rect 439648 37204 439654 37256
rect 132218 35912 132224 35964
rect 132276 35952 132282 35964
rect 186314 35952 186320 35964
rect 132276 35924 186320 35952
rect 132276 35912 132282 35924
rect 186314 35912 186320 35924
rect 186372 35912 186378 35964
rect 131206 35844 131212 35896
rect 131264 35884 131270 35896
rect 186958 35884 186964 35896
rect 131264 35856 186964 35884
rect 131264 35844 131270 35856
rect 186958 35844 186964 35856
rect 187016 35844 187022 35896
rect 417418 35844 417424 35896
rect 417476 35884 417482 35896
rect 437474 35884 437480 35896
rect 417476 35856 437480 35884
rect 417476 35844 417482 35856
rect 437474 35844 437480 35856
rect 437532 35844 437538 35896
rect 131114 35776 131120 35828
rect 131172 35816 131178 35828
rect 187050 35816 187056 35828
rect 131172 35788 187056 35816
rect 131172 35776 131178 35788
rect 187050 35776 187056 35788
rect 187108 35776 187114 35828
rect 411254 35776 411260 35828
rect 411312 35816 411318 35828
rect 418798 35816 418804 35828
rect 411312 35788 418804 35816
rect 411312 35776 411318 35788
rect 418798 35776 418804 35788
rect 418856 35776 418862 35828
rect 414934 34416 414940 34468
rect 414992 34456 414998 34468
rect 437474 34456 437480 34468
rect 414992 34428 437480 34456
rect 414992 34416 414998 34428
rect 437474 34416 437480 34428
rect 437532 34416 437538 34468
rect 131114 33124 131120 33176
rect 131172 33164 131178 33176
rect 186314 33164 186320 33176
rect 131172 33136 186320 33164
rect 131172 33124 131178 33136
rect 186314 33124 186320 33136
rect 186372 33124 186378 33176
rect 131206 33056 131212 33108
rect 131264 33096 131270 33108
rect 186406 33096 186412 33108
rect 131264 33068 186412 33096
rect 131264 33056 131270 33068
rect 186406 33056 186412 33068
rect 186464 33056 186470 33108
rect 412082 33056 412088 33108
rect 412140 33096 412146 33108
rect 437474 33096 437480 33108
rect 412140 33068 437480 33096
rect 412140 33056 412146 33068
rect 437474 33056 437480 33068
rect 437532 33056 437538 33108
rect 411254 32988 411260 33040
rect 411312 33028 411318 33040
rect 418890 33028 418896 33040
rect 411312 33000 418896 33028
rect 411312 32988 411318 33000
rect 418890 32988 418896 33000
rect 418948 32988 418954 33040
rect 131206 31832 131212 31884
rect 131264 31872 131270 31884
rect 186406 31872 186412 31884
rect 131264 31844 186412 31872
rect 131264 31832 131270 31844
rect 186406 31832 186412 31844
rect 186464 31832 186470 31884
rect 131298 31764 131304 31816
rect 131356 31804 131362 31816
rect 186314 31804 186320 31816
rect 131356 31776 186320 31804
rect 131356 31764 131362 31776
rect 186314 31764 186320 31776
rect 186372 31764 186378 31816
rect 411806 31696 411812 31748
rect 411864 31736 411870 31748
rect 542722 31736 542728 31748
rect 411864 31708 542728 31736
rect 411864 31696 411870 31708
rect 542722 31696 542728 31708
rect 542780 31696 542786 31748
rect 412266 31628 412272 31680
rect 412324 31668 412330 31680
rect 542538 31668 542544 31680
rect 412324 31640 542544 31668
rect 412324 31628 412330 31640
rect 542538 31628 542544 31640
rect 542596 31628 542602 31680
rect 412358 31560 412364 31612
rect 412416 31600 412422 31612
rect 542630 31600 542636 31612
rect 412416 31572 542636 31600
rect 412416 31560 412422 31572
rect 542630 31560 542636 31572
rect 542688 31560 542694 31612
rect 412174 31492 412180 31544
rect 412232 31532 412238 31544
rect 437474 31532 437480 31544
rect 412232 31504 437480 31532
rect 412232 31492 412238 31504
rect 437474 31492 437480 31504
rect 437532 31492 437538 31544
rect 131114 31016 131120 31068
rect 131172 31056 131178 31068
rect 186314 31056 186320 31068
rect 131172 31028 186320 31056
rect 131172 31016 131178 31028
rect 186314 31016 186320 31028
rect 186372 31016 186378 31068
rect 439774 30268 439780 30320
rect 439832 30308 439838 30320
rect 542446 30308 542452 30320
rect 439832 30280 542452 30308
rect 439832 30268 439838 30280
rect 542446 30268 542452 30280
rect 542504 30268 542510 30320
rect 439866 30200 439872 30252
rect 439924 30240 439930 30252
rect 542354 30240 542360 30252
rect 439924 30212 542360 30240
rect 439924 30200 439930 30212
rect 542354 30200 542360 30212
rect 542412 30200 542418 30252
rect 131758 29248 131764 29300
rect 131816 29288 131822 29300
rect 283006 29288 283012 29300
rect 131816 29260 283012 29288
rect 131816 29248 131822 29260
rect 283006 29248 283012 29260
rect 283064 29248 283070 29300
rect 440050 29248 440056 29300
rect 440108 29288 440114 29300
rect 484578 29288 484584 29300
rect 440108 29260 484584 29288
rect 440108 29248 440114 29260
rect 484578 29248 484584 29260
rect 484636 29248 484642 29300
rect 130378 29180 130384 29232
rect 130436 29220 130442 29232
rect 316218 29220 316224 29232
rect 130436 29192 316224 29220
rect 130436 29180 130442 29192
rect 316218 29180 316224 29192
rect 316276 29180 316282 29232
rect 438210 29180 438216 29232
rect 438268 29220 438274 29232
rect 524598 29220 524604 29232
rect 438268 29192 524604 29220
rect 438268 29180 438274 29192
rect 524598 29180 524604 29192
rect 524656 29180 524662 29232
rect 206278 29112 206284 29164
rect 206336 29152 206342 29164
rect 410518 29152 410524 29164
rect 206336 29124 410524 29152
rect 206336 29112 206342 29124
rect 410518 29112 410524 29124
rect 410576 29112 410582 29164
rect 435358 29112 435364 29164
rect 435416 29152 435422 29164
rect 534626 29152 534632 29164
rect 435416 29124 534632 29152
rect 435416 29112 435422 29124
rect 534626 29112 534632 29124
rect 534684 29112 534690 29164
rect 130470 29044 130476 29096
rect 130528 29084 130534 29096
rect 371234 29084 371240 29096
rect 130528 29056 371240 29084
rect 130528 29044 130534 29056
rect 371234 29044 371240 29056
rect 371292 29044 371298 29096
rect 413554 29044 413560 29096
rect 413612 29084 413618 29096
rect 514754 29084 514760 29096
rect 413612 29056 514760 29084
rect 413612 29044 413618 29056
rect 514754 29044 514760 29056
rect 514812 29044 514818 29096
rect 205634 28976 205640 29028
rect 205692 29016 205698 29028
rect 206278 29016 206284 29028
rect 205692 28988 206284 29016
rect 205692 28976 205698 28988
rect 206278 28976 206284 28988
rect 206336 28976 206342 29028
rect 217778 28976 217784 29028
rect 217836 29016 217842 29028
rect 540330 29016 540336 29028
rect 217836 28988 540336 29016
rect 217836 28976 217842 28988
rect 540330 28976 540336 28988
rect 540388 28976 540394 29028
rect 79962 28908 79968 28960
rect 80020 28948 80026 28960
rect 464614 28948 464620 28960
rect 80020 28920 464620 28948
rect 80020 28908 80026 28920
rect 464614 28908 464620 28920
rect 464672 28908 464678 28960
rect 195238 28840 195244 28892
rect 195296 28880 195302 28892
rect 439498 28880 439504 28892
rect 195296 28852 439504 28880
rect 195296 28840 195302 28852
rect 439498 28840 439504 28852
rect 439556 28840 439562 28892
rect 445294 28840 445300 28892
rect 445352 28880 445358 28892
rect 540422 28880 540428 28892
rect 445352 28852 540428 28880
rect 445352 28840 445358 28852
rect 540422 28840 540428 28852
rect 540480 28840 540486 28892
rect 188522 28772 188528 28824
rect 188580 28812 188586 28824
rect 404446 28812 404452 28824
rect 188580 28784 404452 28812
rect 188580 28772 188586 28784
rect 404446 28772 404452 28784
rect 404504 28772 404510 28824
rect 413462 28772 413468 28824
rect 413520 28812 413526 28824
rect 504634 28812 504640 28824
rect 413520 28784 504640 28812
rect 413520 28772 413526 28784
rect 504634 28772 504640 28784
rect 504692 28772 504698 28824
rect 188430 28704 188436 28756
rect 188488 28744 188494 28756
rect 393406 28744 393412 28756
rect 188488 28716 393412 28744
rect 188488 28704 188494 28716
rect 393406 28704 393412 28716
rect 393464 28704 393470 28756
rect 455230 28704 455236 28756
rect 455288 28744 455294 28756
rect 541618 28744 541624 28756
rect 455288 28716 541624 28744
rect 455288 28704 455294 28716
rect 541618 28704 541624 28716
rect 541676 28704 541682 28756
rect 166258 28636 166264 28688
rect 166316 28676 166322 28688
rect 360194 28676 360200 28688
rect 166316 28648 360200 28676
rect 166316 28636 166322 28648
rect 360194 28636 360200 28648
rect 360252 28636 360258 28688
rect 411254 28636 411260 28688
rect 411312 28676 411318 28688
rect 474734 28676 474740 28688
rect 411312 28648 474740 28676
rect 411312 28636 411318 28648
rect 474734 28636 474740 28648
rect 474792 28636 474798 28688
rect 189994 28568 190000 28620
rect 190052 28608 190058 28620
rect 382274 28608 382280 28620
rect 190052 28580 382280 28608
rect 190052 28568 190058 28580
rect 382274 28568 382280 28580
rect 382332 28568 382338 28620
rect 439958 28568 439964 28620
rect 440016 28608 440022 28620
rect 494606 28608 494612 28620
rect 440016 28580 494612 28608
rect 440016 28568 440022 28580
rect 494606 28568 494612 28580
rect 494664 28568 494670 28620
rect 164878 28500 164884 28552
rect 164936 28540 164942 28552
rect 349154 28540 349160 28552
rect 164936 28512 349160 28540
rect 164936 28500 164942 28512
rect 349154 28500 349160 28512
rect 349212 28500 349218 28552
rect 188338 28432 188344 28484
rect 188396 28472 188402 28484
rect 338114 28472 338120 28484
rect 188396 28444 338120 28472
rect 188396 28432 188402 28444
rect 338114 28432 338120 28444
rect 338172 28432 338178 28484
rect 189902 28364 189908 28416
rect 189960 28404 189966 28416
rect 327074 28404 327080 28416
rect 189960 28376 327080 28404
rect 189960 28364 189966 28376
rect 327074 28364 327080 28376
rect 327132 28364 327138 28416
rect 133138 28296 133144 28348
rect 133196 28336 133202 28348
rect 239030 28336 239036 28348
rect 133196 28308 239036 28336
rect 133196 28296 133202 28308
rect 239030 28296 239036 28308
rect 239088 28296 239094 28348
rect 190086 28228 190092 28280
rect 190144 28268 190150 28280
rect 294046 28268 294052 28280
rect 190144 28240 294052 28268
rect 190144 28228 190150 28240
rect 294046 28228 294052 28240
rect 294104 28228 294110 28280
rect 189718 28160 189724 28212
rect 189776 28200 189782 28212
rect 271966 28200 271972 28212
rect 189776 28172 271972 28200
rect 189776 28160 189782 28172
rect 271966 28160 271972 28172
rect 272024 28160 272030 28212
rect 189810 28092 189816 28144
rect 189868 28132 189874 28144
rect 261110 28132 261116 28144
rect 189868 28104 261116 28132
rect 189868 28092 189874 28104
rect 261110 28092 261116 28104
rect 261168 28092 261174 28144
rect 190178 28024 190184 28076
rect 190236 28064 190242 28076
rect 250070 28064 250076 28076
rect 190236 28036 250076 28064
rect 190236 28024 190242 28036
rect 250070 28024 250076 28036
rect 250128 28024 250134 28076
rect 540238 20612 540244 20664
rect 540296 20652 540302 20664
rect 579982 20652 579988 20664
rect 540296 20624 579988 20652
rect 540296 20612 540302 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 227714 6808 227720 6860
rect 227772 6848 227778 6860
rect 580166 6848 580172 6860
rect 227772 6820 580172 6848
rect 227772 6808 227778 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 2682 4088 2688 4140
rect 2740 4128 2746 4140
rect 205634 4128 205640 4140
rect 2740 4100 205640 4128
rect 2740 4088 2746 4100
rect 205634 4088 205640 4100
rect 205692 4088 205698 4140
rect 1302 4020 1308 4072
rect 1360 4060 1366 4072
rect 195238 4060 195244 4072
rect 1360 4032 195244 4060
rect 1360 4020 1366 4032
rect 195238 4020 195244 4032
rect 195296 4020 195302 4072
rect 1670 3680 1676 3732
rect 1728 3720 1734 3732
rect 2682 3720 2688 3732
rect 1728 3692 2688 3720
rect 1728 3680 1734 3692
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 566 3612 572 3664
rect 624 3652 630 3664
rect 1302 3652 1308 3664
rect 624 3624 1308 3652
rect 624 3612 630 3624
rect 1302 3612 1308 3624
rect 1360 3612 1366 3664
<< via1 >>
rect 204260 325660 204312 325712
rect 207020 325660 207072 325712
rect 193220 306348 193272 306400
rect 207020 306348 207072 306400
rect 190460 304988 190512 305040
rect 207020 304988 207072 305040
rect 67824 298256 67876 298308
rect 227720 298256 227772 298308
rect 69296 298188 69348 298240
rect 229100 298188 229152 298240
rect 55220 298120 55272 298172
rect 55864 298120 55916 298172
rect 215852 298120 215904 298172
rect 76840 297984 76892 298036
rect 79324 297984 79376 298036
rect 97080 297440 97132 297492
rect 130476 297440 130528 297492
rect 89168 297372 89220 297424
rect 130384 297372 130436 297424
rect 75552 297304 75604 297356
rect 131764 297304 131816 297356
rect 70216 297236 70268 297288
rect 229284 297236 229336 297288
rect 106648 297168 106700 297220
rect 341524 297168 341576 297220
rect 107752 297100 107804 297152
rect 345664 297100 345716 297152
rect 111616 297032 111668 297084
rect 409052 297032 409104 297084
rect 105544 296964 105596 297016
rect 408868 296964 408920 297016
rect 104256 296896 104308 296948
rect 409328 296896 409380 296948
rect 102968 296828 103020 296880
rect 409236 296828 409288 296880
rect 102048 296760 102100 296812
rect 409144 296760 409196 296812
rect 65800 296692 65852 296744
rect 408960 296692 409012 296744
rect 234620 295944 234672 295996
rect 242900 295944 242952 295996
rect 49424 291796 49476 291848
rect 371240 291796 371292 291848
rect 47768 287648 47820 287700
rect 409972 287648 410024 287700
rect 208124 282344 208176 282396
rect 213920 282344 213972 282396
rect 194600 282276 194652 282328
rect 224960 282276 225012 282328
rect 266176 282276 266228 282328
rect 358820 282276 358872 282328
rect 197360 282208 197412 282260
rect 237380 282208 237432 282260
rect 267464 282208 267516 282260
rect 364340 282208 364392 282260
rect 47860 282140 47912 282192
rect 410064 282140 410116 282192
rect 218060 280848 218112 280900
rect 229100 280848 229152 280900
rect 209596 280780 209648 280832
rect 231860 280780 231912 280832
rect 248236 280780 248288 280832
rect 259460 280780 259512 280832
rect 209504 279624 209556 279676
rect 222200 279624 222252 279676
rect 85304 279556 85356 279608
rect 389180 279556 389232 279608
rect 49516 279488 49568 279540
rect 374000 279488 374052 279540
rect 47676 279420 47728 279472
rect 409880 279420 409932 279472
rect 245568 273912 245620 273964
rect 280160 273912 280212 273964
rect 246764 271804 246816 271856
rect 248420 271804 248472 271856
rect 264796 268404 264848 268456
rect 354680 268404 354732 268456
rect 242808 268336 242860 268388
rect 266360 268336 266412 268388
rect 267556 268336 267608 268388
rect 368480 268336 368532 268388
rect 229100 268132 229152 268184
rect 234712 268132 234764 268184
rect 260656 267112 260708 267164
rect 341064 267112 341116 267164
rect 262036 267044 262088 267096
rect 345572 267044 345624 267096
rect 263416 266976 263468 267028
rect 350540 266976 350592 267028
rect 257804 265752 257856 265804
rect 327264 265752 327316 265804
rect 259276 265684 259328 265736
rect 331864 265684 331916 265736
rect 259184 265616 259236 265668
rect 336740 265616 336792 265668
rect 253756 264392 253808 264444
rect 313280 264392 313332 264444
rect 255136 264324 255188 264376
rect 318064 264324 318116 264376
rect 256516 264256 256568 264308
rect 322940 264256 322992 264308
rect 100576 264188 100628 264240
rect 399024 264188 399076 264240
rect 248328 263100 248380 263152
rect 290280 263100 290332 263152
rect 252284 263032 252336 263084
rect 304080 263032 304132 263084
rect 252376 262964 252428 263016
rect 309232 262964 309284 263016
rect 96436 262896 96488 262948
rect 411904 262896 411956 262948
rect 81256 262828 81308 262880
rect 411536 262828 411588 262880
rect 255228 261808 255280 261860
rect 283288 261808 283340 261860
rect 256608 261740 256660 261792
rect 287888 261740 287940 261792
rect 211528 261672 211580 261724
rect 231952 261672 232004 261724
rect 246856 261672 246908 261724
rect 255504 261672 255556 261724
rect 259368 261672 259420 261724
rect 302332 261672 302384 261724
rect 88156 261604 88208 261656
rect 387800 261604 387852 261656
rect 90916 261536 90968 261588
rect 392032 261536 392084 261588
rect 86684 261468 86736 261520
rect 411628 261468 411680 261520
rect 252468 260448 252520 260500
rect 274088 260448 274140 260500
rect 225328 260380 225380 260432
rect 241520 260380 241572 260432
rect 253848 260380 253900 260432
rect 278780 260380 278832 260432
rect 74448 260312 74500 260364
rect 148324 260312 148376 260364
rect 216128 260312 216180 260364
rect 240140 260312 240192 260364
rect 273076 260312 273128 260364
rect 348056 260312 348108 260364
rect 79876 260244 79928 260296
rect 153200 260244 153252 260296
rect 202144 260244 202196 260296
rect 230480 260244 230532 260296
rect 237196 260244 237248 260296
rect 244372 260244 244424 260296
rect 250996 260244 251048 260296
rect 269304 260244 269356 260296
rect 273168 260244 273220 260296
rect 352656 260244 352708 260296
rect 115848 260176 115900 260228
rect 403624 260176 403676 260228
rect 112996 260108 113048 260160
rect 401600 260108 401652 260160
rect 241612 260040 241664 260092
rect 244280 260040 244332 260092
rect 244096 258952 244148 259004
rect 276296 258952 276348 259004
rect 249616 258884 249668 258936
rect 294880 258884 294932 258936
rect 251088 258816 251140 258868
rect 299480 258816 299532 258868
rect 93584 258748 93636 258800
rect 410248 258748 410300 258800
rect 85396 258680 85448 258732
rect 411352 258680 411404 258732
rect 246948 257660 247000 257712
rect 285680 257660 285732 257712
rect 260748 257592 260800 257644
rect 306564 257592 306616 257644
rect 244188 257524 244240 257576
rect 271880 257524 271932 257576
rect 277308 257524 277360 257576
rect 366732 257524 366784 257576
rect 108856 257456 108908 257508
rect 396724 257456 396776 257508
rect 104716 257388 104768 257440
rect 394700 257388 394752 257440
rect 81348 257320 81400 257372
rect 375932 257320 375984 257372
rect 221464 256232 221516 256284
rect 233240 256232 233292 256284
rect 257896 256232 257948 256284
rect 297180 256232 297232 256284
rect 209504 256164 209556 256216
rect 227720 256164 227772 256216
rect 262128 256164 262180 256216
rect 311164 256164 311216 256216
rect 201408 256096 201460 256148
rect 226340 256096 226392 256148
rect 263508 256096 263560 256148
rect 316040 256096 316092 256148
rect 97816 256028 97868 256080
rect 410432 256028 410484 256080
rect 84016 255960 84068 256012
rect 411444 255960 411496 256012
rect 209688 254736 209740 254788
rect 253204 254736 253256 254788
rect 257988 254736 258040 254788
rect 292580 254736 292632 254788
rect 92296 254668 92348 254720
rect 410340 254668 410392 254720
rect 91008 254600 91060 254652
rect 410156 254600 410208 254652
rect 82636 254532 82688 254584
rect 411260 254532 411312 254584
rect 228456 253852 228508 253904
rect 229192 253852 229244 253904
rect 264888 253648 264940 253700
rect 320364 253648 320416 253700
rect 266268 253580 266320 253632
rect 324964 253580 325016 253632
rect 267648 253512 267700 253564
rect 329840 253512 329892 253564
rect 269028 253444 269080 253496
rect 334348 253444 334400 253496
rect 208216 253376 208268 253428
rect 239404 253376 239456 253428
rect 270408 253376 270460 253428
rect 338948 253376 339000 253428
rect 271788 253308 271840 253360
rect 343640 253308 343692 253360
rect 207664 253240 207716 253292
rect 238760 253240 238812 253292
rect 240048 253240 240100 253292
rect 258080 253240 258132 253292
rect 274548 253240 274600 253292
rect 357532 253240 357584 253292
rect 208308 253172 208360 253224
rect 246396 253172 246448 253224
rect 249708 253172 249760 253224
rect 264980 253172 265032 253224
rect 275928 253172 275980 253224
rect 362132 253172 362184 253224
rect 67548 252492 67600 252544
rect 200396 252492 200448 252544
rect 201408 252492 201460 252544
rect 238668 252152 238720 252204
rect 251180 252152 251232 252204
rect 345664 252152 345716 252204
rect 408500 252152 408552 252204
rect 241428 252084 241480 252136
rect 262588 252084 262640 252136
rect 341524 252084 341576 252136
rect 406108 252084 406160 252136
rect 148324 252016 148376 252068
rect 378324 252016 378376 252068
rect 153200 251948 153252 252000
rect 385316 251948 385368 252000
rect 79324 251880 79376 251932
rect 380992 251880 381044 251932
rect 77116 251812 77168 251864
rect 382924 251812 382976 251864
rect 101956 250588 102008 250640
rect 410524 250588 410576 250640
rect 82728 250520 82780 250572
rect 411812 250520 411864 250572
rect 78496 250452 78548 250504
rect 411720 250452 411772 250504
rect 114468 249704 114520 249756
rect 186320 249704 186372 249756
rect 106096 248344 106148 248396
rect 186412 248344 186464 248396
rect 107476 248276 107528 248328
rect 186320 248276 186372 248328
rect 95056 246984 95108 247036
rect 186320 246984 186372 247036
rect 85488 246304 85540 246356
rect 187148 246304 187200 246356
rect 103336 245556 103388 245608
rect 186320 245556 186372 245608
rect 101864 244196 101916 244248
rect 186320 244196 186372 244248
rect 100668 242836 100720 242888
rect 186320 242836 186372 242888
rect 88248 241408 88300 241460
rect 186320 241408 186372 241460
rect 95148 240048 95200 240100
rect 186412 240048 186464 240100
rect 96528 239980 96580 240032
rect 186320 239980 186372 240032
rect 84108 237328 84160 237380
rect 186320 237328 186372 237380
rect 89536 235900 89588 235952
rect 186320 235900 186372 235952
rect 86776 234540 86828 234592
rect 186320 234540 186372 234592
rect 49608 233180 49660 233232
rect 186412 233180 186464 233232
rect 86868 233112 86920 233164
rect 186320 233112 186372 233164
rect 73068 231752 73120 231804
rect 186320 231752 186372 231804
rect 71688 230392 71740 230444
rect 186320 230392 186372 230444
rect 169024 227740 169076 227792
rect 186320 227740 186372 227792
rect 148324 226312 148376 226364
rect 186320 226312 186372 226364
rect 157984 225020 158036 225072
rect 186412 225020 186464 225072
rect 133236 224952 133288 225004
rect 186320 224952 186372 225004
rect 151084 223592 151136 223644
rect 186320 223592 186372 223644
rect 145564 222164 145616 222216
rect 186320 222164 186372 222216
rect 162124 220804 162176 220856
rect 186320 220804 186372 220856
rect 145656 219444 145708 219496
rect 186320 219444 186372 219496
rect 156604 218084 156656 218136
rect 186412 218084 186464 218136
rect 135904 218016 135956 218068
rect 186320 218016 186372 218068
rect 543004 218016 543056 218068
rect 580172 218016 580224 218068
rect 149704 216656 149756 216708
rect 186320 216656 186372 216708
rect 142804 215296 142856 215348
rect 186320 215296 186372 215348
rect 155224 213936 155276 213988
rect 186320 213936 186372 213988
rect 135996 212508 136048 212560
rect 186320 212508 186372 212560
rect 145748 211148 145800 211200
rect 186320 211148 186372 211200
rect 160744 209856 160796 209908
rect 186320 209856 186372 209908
rect 149796 209788 149848 209840
rect 186412 209788 186464 209840
rect 159364 207000 159416 207052
rect 186320 207000 186372 207052
rect 158076 205640 158128 205692
rect 186320 205640 186372 205692
rect 140044 204280 140096 204332
rect 186320 204280 186372 204332
rect 146944 202920 146996 202972
rect 186320 202920 186372 202972
rect 134616 202852 134668 202904
rect 186412 202852 186464 202904
rect 411260 202852 411312 202904
rect 540244 202852 540296 202904
rect 411260 201560 411312 201612
rect 414664 201560 414716 201612
rect 134524 201492 134576 201544
rect 186320 201492 186372 201544
rect 144184 200132 144236 200184
rect 186320 200132 186372 200184
rect 134708 198704 134760 198756
rect 186320 198704 186372 198756
rect 411260 198704 411312 198756
rect 540336 198704 540388 198756
rect 159456 197344 159508 197396
rect 186320 197344 186372 197396
rect 411260 197344 411312 197396
rect 540428 197344 540480 197396
rect 147036 194624 147088 194676
rect 186320 194624 186372 194676
rect 141424 194556 141476 194608
rect 186412 194556 186464 194608
rect 411260 193536 411312 193588
rect 413376 193536 413428 193588
rect 137284 193196 137336 193248
rect 186320 193196 186372 193248
rect 147128 191836 147180 191888
rect 186320 191836 186372 191888
rect 93676 191224 93728 191276
rect 166264 191224 166316 191276
rect 92388 191156 92440 191208
rect 188344 191156 188396 191208
rect 79968 191088 80020 191140
rect 189724 191088 189776 191140
rect 140136 190476 140188 190528
rect 186320 190476 186372 190528
rect 156696 189048 156748 189100
rect 186320 189048 186372 189100
rect 411260 189048 411312 189100
rect 428464 189048 428516 189100
rect 159548 187756 159600 187808
rect 186412 187756 186464 187808
rect 133328 187688 133380 187740
rect 186320 187688 186372 187740
rect 411260 187688 411312 187740
rect 428556 187688 428608 187740
rect 137376 186328 137428 186380
rect 186320 186328 186372 186380
rect 411260 186328 411312 186380
rect 418988 186328 419040 186380
rect 141516 184900 141568 184952
rect 186320 184900 186372 184952
rect 140228 183540 140280 183592
rect 186320 183540 186372 183592
rect 411260 183540 411312 183592
rect 428648 183540 428700 183592
rect 156880 182180 156932 182232
rect 186320 182180 186372 182232
rect 411260 182180 411312 182232
rect 436744 182180 436796 182232
rect 156788 180888 156840 180940
rect 186320 180888 186372 180940
rect 140320 180820 140372 180872
rect 186412 180820 186464 180872
rect 137468 179392 137520 179444
rect 186320 179392 186372 179444
rect 411260 179392 411312 179444
rect 425704 179392 425756 179444
rect 144276 178032 144328 178084
rect 186320 178032 186372 178084
rect 411260 178032 411312 178084
rect 435364 178032 435416 178084
rect 543096 178032 543148 178084
rect 580172 178032 580224 178084
rect 138664 176672 138716 176724
rect 186320 176672 186372 176724
rect 411260 176672 411312 176724
rect 417424 176672 417476 176724
rect 141608 175244 141660 175296
rect 186320 175244 186372 175296
rect 411260 174428 411312 174480
rect 414940 174428 414992 174480
rect 164976 173884 165028 173936
rect 186320 173884 186372 173936
rect 160836 172592 160888 172644
rect 186320 172592 186372 172644
rect 138756 172524 138808 172576
rect 186412 172524 186464 172576
rect 411260 172524 411312 172576
rect 432604 172524 432656 172576
rect 137560 171096 137612 171148
rect 186320 171096 186372 171148
rect 411260 171096 411312 171148
rect 431224 171096 431276 171148
rect 131856 169736 131908 169788
rect 186320 169736 186372 169788
rect 158168 168376 158220 168428
rect 186320 168376 186372 168428
rect 411260 168376 411312 168428
rect 429844 168376 429896 168428
rect 162216 167016 162268 167068
rect 186320 167016 186372 167068
rect 411260 167016 411312 167068
rect 428740 167016 428792 167068
rect 159640 165656 159692 165708
rect 186320 165656 186372 165708
rect 158260 165588 158312 165640
rect 186412 165588 186464 165640
rect 155316 164228 155368 164280
rect 186320 164228 186372 164280
rect 411260 164228 411312 164280
rect 425796 164228 425848 164280
rect 160928 162868 160980 162920
rect 186320 162868 186372 162920
rect 411260 162868 411312 162920
rect 424324 162868 424376 162920
rect 134800 161440 134852 161492
rect 186320 161440 186372 161492
rect 411260 161440 411312 161492
rect 424416 161440 424468 161492
rect 158352 160080 158404 160132
rect 186320 160080 186372 160132
rect 133512 158720 133564 158772
rect 186320 158720 186372 158772
rect 411260 158720 411312 158772
rect 423128 158720 423180 158772
rect 156972 157428 157024 157480
rect 186412 157428 186464 157480
rect 133420 157360 133472 157412
rect 186320 157360 186372 157412
rect 411260 157360 411312 157412
rect 425888 157360 425940 157412
rect 136088 155932 136140 155984
rect 186320 155932 186372 155984
rect 411260 155932 411312 155984
rect 423036 155932 423088 155984
rect 133604 154572 133656 154624
rect 186320 154572 186372 154624
rect 138848 153212 138900 153264
rect 186320 153212 186372 153264
rect 411260 153212 411312 153264
rect 417516 153212 417568 153264
rect 141700 151784 141752 151836
rect 186320 151784 186372 151836
rect 411260 151784 411312 151836
rect 422944 151784 422996 151836
rect 166356 150492 166408 150544
rect 186412 150492 186464 150544
rect 155408 150424 155460 150476
rect 186320 150424 186372 150476
rect 151176 149064 151228 149116
rect 186320 149064 186372 149116
rect 411260 149064 411312 149116
rect 417608 149064 417660 149116
rect 144368 147636 144420 147688
rect 186320 147636 186372 147688
rect 411260 147636 411312 147688
rect 421656 147636 421708 147688
rect 155500 146276 155552 146328
rect 186320 146276 186372 146328
rect 411260 146276 411312 146328
rect 419172 146276 419224 146328
rect 151268 144916 151320 144968
rect 186320 144916 186372 144968
rect 152464 143624 152516 143676
rect 186320 143624 186372 143676
rect 144460 143556 144512 143608
rect 186412 143556 186464 143608
rect 411260 143556 411312 143608
rect 421564 143556 421616 143608
rect 148416 142128 148468 142180
rect 186320 142128 186372 142180
rect 411260 142128 411312 142180
rect 429936 142128 429988 142180
rect 411260 140768 411312 140820
rect 417700 140768 417752 140820
rect 152556 139408 152608 139460
rect 186320 139408 186372 139460
rect 414664 139340 414716 139392
rect 580172 139340 580224 139392
rect 148508 137980 148560 138032
rect 186320 137980 186372 138032
rect 411260 137980 411312 138032
rect 426072 137980 426124 138032
rect 142896 136620 142948 136672
rect 186320 136620 186372 136672
rect 411260 136620 411312 136672
rect 425980 136620 426032 136672
rect 152648 135328 152700 135380
rect 186412 135328 186464 135380
rect 148600 135260 148652 135312
rect 186320 135260 186372 135312
rect 411260 135260 411312 135312
rect 431316 135260 431368 135312
rect 93768 133288 93820 133340
rect 164884 133288 164936 133340
rect 117228 133220 117280 133272
rect 188528 133220 188580 133272
rect 113088 133152 113140 133204
rect 188436 133152 188488 133204
rect 152740 132472 152792 132524
rect 186320 132472 186372 132524
rect 411260 132472 411312 132524
rect 424508 132472 424560 132524
rect 110328 131860 110380 131912
rect 190000 131860 190052 131912
rect 97908 131792 97960 131844
rect 189908 131792 189960 131844
rect 48136 131724 48188 131776
rect 189816 131724 189868 131776
rect 413468 131452 413520 131504
rect 521752 131452 521804 131504
rect 439688 131384 439740 131436
rect 472072 131384 472124 131436
rect 414664 131316 414716 131368
rect 478880 131316 478932 131368
rect 414756 131248 414808 131300
rect 485964 131248 486016 131300
rect 1308 131180 1360 131232
rect 55128 131180 55180 131232
rect 438124 131180 438176 131232
rect 536012 131180 536064 131232
rect 2688 131112 2740 131164
rect 104900 131112 104952 131164
rect 148692 131112 148744 131164
rect 186320 131112 186372 131164
rect 411260 131112 411312 131164
rect 415032 131112 415084 131164
rect 439504 131112 439556 131164
rect 443184 131112 443236 131164
rect 48044 130500 48096 130552
rect 133144 130500 133196 130552
rect 78588 130432 78640 130484
rect 190184 130432 190236 130484
rect 439872 130432 439924 130484
rect 542544 130432 542596 130484
rect 48228 130364 48280 130416
rect 190092 130364 190144 130416
rect 438768 130364 438820 130416
rect 450268 130364 450320 130416
rect 439596 130296 439648 130348
rect 464528 130296 464580 130348
rect 419080 130228 419132 130280
rect 493140 130228 493192 130280
rect 439780 130160 439832 130212
rect 514898 130160 514950 130212
rect 420184 130092 420236 130144
rect 500638 130092 500690 130144
rect 420276 130024 420328 130076
rect 507400 130024 507452 130076
rect 435548 129956 435600 130008
rect 528836 129956 528888 130008
rect 439964 129888 440016 129940
rect 539324 129888 539376 129940
rect 418804 129820 418856 129872
rect 457444 129820 457496 129872
rect 142988 129752 143040 129804
rect 186320 129752 186372 129804
rect 412272 129752 412324 129804
rect 542360 129752 542412 129804
rect 131120 129684 131172 129736
rect 169024 129684 169076 129736
rect 131304 129616 131356 129668
rect 157984 129616 158036 129668
rect 131212 129548 131264 129600
rect 148324 129548 148376 129600
rect 411260 128460 411312 128512
rect 424600 128460 424652 128512
rect 151360 128392 151412 128444
rect 186412 128392 186464 128444
rect 421932 128392 421984 128444
rect 437480 128392 437532 128444
rect 147220 128324 147272 128376
rect 186320 128324 186372 128376
rect 412364 128324 412416 128376
rect 542452 128324 542504 128376
rect 132040 128256 132092 128308
rect 151084 128256 151136 128308
rect 132224 128188 132276 128240
rect 133236 128188 133288 128240
rect 411260 127032 411312 127084
rect 432696 127032 432748 127084
rect 143080 126964 143132 127016
rect 186320 126964 186372 127016
rect 413560 126964 413612 127016
rect 437480 126964 437532 127016
rect 131120 126896 131172 126948
rect 162124 126896 162176 126948
rect 132040 126828 132092 126880
rect 145656 126828 145708 126880
rect 131212 126760 131264 126812
rect 145564 126760 145616 126812
rect 411260 125672 411312 125724
rect 416044 125672 416096 125724
rect 151084 125604 151136 125656
rect 186320 125604 186372 125656
rect 413652 125604 413704 125656
rect 437480 125604 437532 125656
rect 541624 125604 541676 125656
rect 580172 125604 580224 125656
rect 131120 125536 131172 125588
rect 156604 125536 156656 125588
rect 131212 125468 131264 125520
rect 135904 125468 135956 125520
rect 436100 124448 436152 124500
rect 438768 124448 438820 124500
rect 145564 124176 145616 124228
rect 186320 124176 186372 124228
rect 414848 124176 414900 124228
rect 437480 124176 437532 124228
rect 132224 124108 132276 124160
rect 149704 124108 149756 124160
rect 131120 124040 131172 124092
rect 142804 124040 142856 124092
rect 411260 122816 411312 122868
rect 435456 122816 435508 122868
rect 131212 122748 131264 122800
rect 155224 122748 155276 122800
rect 131120 122680 131172 122732
rect 145748 122680 145800 122732
rect 131212 122612 131264 122664
rect 135996 122612 136048 122664
rect 411260 121524 411312 121576
rect 416136 121524 416188 121576
rect 149704 121456 149756 121508
rect 186320 121456 186372 121508
rect 413284 121456 413336 121508
rect 437480 121456 437532 121508
rect 131948 121388 132000 121440
rect 160744 121388 160796 121440
rect 131212 121320 131264 121372
rect 149796 121320 149848 121372
rect 145748 120164 145800 120216
rect 186412 120164 186464 120216
rect 434076 120164 434128 120216
rect 436008 120164 436060 120216
rect 142804 120096 142856 120148
rect 186320 120096 186372 120148
rect 418896 120096 418948 120148
rect 437480 120096 437532 120148
rect 132224 120028 132276 120080
rect 186964 120028 187016 120080
rect 411996 120028 412048 120080
rect 437572 120028 437624 120080
rect 131120 119960 131172 120012
rect 159364 119960 159416 120012
rect 135904 118668 135956 118720
rect 186320 118668 186372 118720
rect 411260 118668 411312 118720
rect 424692 118668 424744 118720
rect 131212 118600 131264 118652
rect 158076 118600 158128 118652
rect 413376 118600 413428 118652
rect 437480 118600 437532 118652
rect 131120 118532 131172 118584
rect 140044 118532 140096 118584
rect 131212 118464 131264 118516
rect 134616 118464 134668 118516
rect 145656 117308 145708 117360
rect 186320 117308 186372 117360
rect 411260 117308 411312 117360
rect 436836 117308 436888 117360
rect 131212 117240 131264 117292
rect 146944 117240 146996 117292
rect 131120 117172 131172 117224
rect 134524 117172 134576 117224
rect 141792 115948 141844 116000
rect 186320 115948 186372 116000
rect 411260 115948 411312 116000
rect 423220 115948 423272 116000
rect 131212 115880 131264 115932
rect 144184 115880 144236 115932
rect 411904 115880 411956 115932
rect 437480 115880 437532 115932
rect 131212 115472 131264 115524
rect 134708 115472 134760 115524
rect 431960 115200 432012 115252
rect 434076 115200 434128 115252
rect 149796 114520 149848 114572
rect 186320 114520 186372 114572
rect 131304 114452 131356 114504
rect 187056 114452 187108 114504
rect 428464 114452 428516 114504
rect 437480 114452 437532 114504
rect 131212 114384 131264 114436
rect 159456 114384 159508 114436
rect 131120 114316 131172 114368
rect 141424 114316 141476 114368
rect 131212 113092 131264 113144
rect 147036 113092 147088 113144
rect 428556 113092 428608 113144
rect 437480 113092 437532 113144
rect 131120 113024 131172 113076
rect 137284 113024 137336 113076
rect 146944 111800 146996 111852
rect 186320 111800 186372 111852
rect 411260 111800 411312 111852
rect 421840 111800 421892 111852
rect 132132 111732 132184 111784
rect 147128 111732 147180 111784
rect 418988 111732 419040 111784
rect 437480 111732 437532 111784
rect 131212 111664 131264 111716
rect 140136 111664 140188 111716
rect 134524 110440 134576 110492
rect 186320 110440 186372 110492
rect 411260 110440 411312 110492
rect 421748 110440 421800 110492
rect 131304 110372 131356 110424
rect 133328 110372 133380 110424
rect 427820 110372 427872 110424
rect 431868 110440 431920 110492
rect 131212 110304 131264 110356
rect 156696 110304 156748 110356
rect 428648 110304 428700 110356
rect 437480 110304 437532 110356
rect 131120 110236 131172 110288
rect 159548 110236 159600 110288
rect 141424 109012 141476 109064
rect 186320 109012 186372 109064
rect 131120 108944 131172 108996
rect 141516 108944 141568 108996
rect 131212 108876 131264 108928
rect 137376 108876 137428 108928
rect 424968 108060 425020 108112
rect 427820 108060 427872 108112
rect 147036 107652 147088 107704
rect 186320 107652 186372 107704
rect 131120 107584 131172 107636
rect 156880 107584 156932 107636
rect 131304 107516 131356 107568
rect 140320 107516 140372 107568
rect 131212 107448 131264 107500
rect 140228 107448 140280 107500
rect 418160 106700 418212 106752
rect 424968 106700 425020 106752
rect 147128 106360 147180 106412
rect 186412 106360 186464 106412
rect 140044 106292 140096 106344
rect 186320 106292 186372 106344
rect 411260 106292 411312 106344
rect 417792 106292 417844 106344
rect 131120 106224 131172 106276
rect 156788 106224 156840 106276
rect 425704 106224 425756 106276
rect 437480 106224 437532 106276
rect 131212 106156 131264 106208
rect 137468 106156 137520 106208
rect 141516 104864 141568 104916
rect 186320 104864 186372 104916
rect 131212 104796 131264 104848
rect 144276 104796 144328 104848
rect 435364 104796 435416 104848
rect 437664 104796 437716 104848
rect 131120 104728 131172 104780
rect 138664 104728 138716 104780
rect 134616 103504 134668 103556
rect 186320 103504 186372 103556
rect 411260 103504 411312 103556
rect 413376 103504 413428 103556
rect 131672 103436 131724 103488
rect 164976 103436 165028 103488
rect 417424 103436 417476 103488
rect 437480 103436 437532 103488
rect 131212 103368 131264 103420
rect 141608 103368 141660 103420
rect 131120 103300 131172 103352
rect 138756 103300 138808 103352
rect 140136 102144 140188 102196
rect 186320 102144 186372 102196
rect 411260 102144 411312 102196
rect 418988 102144 419040 102196
rect 131212 102076 131264 102128
rect 160836 102076 160888 102128
rect 414940 102076 414992 102128
rect 437480 102076 437532 102128
rect 131120 102008 131172 102060
rect 137560 102008 137612 102060
rect 133696 101396 133748 101448
rect 187424 101396 187476 101448
rect 134708 100716 134760 100768
rect 186320 100716 186372 100768
rect 411260 100716 411312 100768
rect 417424 100716 417476 100768
rect 131212 100648 131264 100700
rect 158168 100648 158220 100700
rect 540428 100648 540480 100700
rect 580172 100648 580224 100700
rect 131488 99968 131540 100020
rect 159640 99968 159692 100020
rect 144184 99356 144236 99408
rect 186320 99356 186372 99408
rect 415952 99356 416004 99408
rect 417884 99356 417936 99408
rect 131212 99288 131264 99340
rect 162216 99288 162268 99340
rect 432604 99288 432656 99340
rect 437480 99288 437532 99340
rect 131120 99220 131172 99272
rect 158260 99220 158312 99272
rect 141608 98064 141660 98116
rect 186412 98064 186464 98116
rect 131856 97996 131908 98048
rect 186320 97996 186372 98048
rect 411260 97996 411312 98048
rect 414940 97996 414992 98048
rect 131120 97928 131172 97980
rect 160928 97928 160980 97980
rect 431224 97928 431276 97980
rect 437480 97928 437532 97980
rect 131212 97860 131264 97912
rect 155316 97860 155368 97912
rect 140228 96636 140280 96688
rect 186320 96636 186372 96688
rect 131120 96568 131172 96620
rect 158352 96568 158404 96620
rect 429844 96568 429896 96620
rect 437480 96568 437532 96620
rect 131212 96432 131264 96484
rect 134800 96432 134852 96484
rect 414020 96024 414072 96076
rect 415952 96024 416004 96076
rect 132224 95956 132276 96008
rect 133512 95956 133564 96008
rect 140320 95208 140372 95260
rect 186320 95208 186372 95260
rect 131212 95140 131264 95192
rect 156972 95140 157024 95192
rect 428740 95140 428792 95192
rect 437480 95140 437532 95192
rect 131120 95072 131172 95124
rect 133420 95072 133472 95124
rect 131948 93848 132000 93900
rect 186320 93848 186372 93900
rect 131212 93780 131264 93832
rect 136088 93780 136140 93832
rect 425796 93780 425848 93832
rect 437480 93780 437532 93832
rect 131120 93712 131172 93764
rect 133604 93712 133656 93764
rect 133236 92488 133288 92540
rect 186320 92488 186372 92540
rect 411352 92488 411404 92540
rect 435364 92488 435416 92540
rect 131304 92420 131356 92472
rect 166356 92420 166408 92472
rect 411260 92420 411312 92472
rect 421932 92420 421984 92472
rect 131120 92352 131172 92404
rect 141700 92352 141752 92404
rect 131212 92284 131264 92336
rect 138848 92284 138900 92336
rect 181444 91060 181496 91112
rect 186320 91060 186372 91112
rect 131212 90992 131264 91044
rect 155408 90992 155460 91044
rect 410524 90992 410576 91044
rect 414020 91060 414072 91112
rect 424324 90992 424376 91044
rect 437480 90992 437532 91044
rect 131120 90924 131172 90976
rect 151176 90924 151228 90976
rect 415032 90312 415084 90364
rect 438308 90312 438360 90364
rect 133328 89700 133380 89752
rect 186320 89700 186372 89752
rect 131304 89632 131356 89684
rect 155500 89632 155552 89684
rect 411260 89632 411312 89684
rect 413560 89632 413612 89684
rect 424416 89632 424468 89684
rect 437480 89632 437532 89684
rect 132224 89564 132276 89616
rect 144368 89564 144420 89616
rect 131120 88952 131172 89004
rect 144460 88952 144512 89004
rect 411812 88952 411864 89004
rect 412180 88952 412232 89004
rect 138664 88340 138716 88392
rect 186320 88340 186372 88392
rect 131304 88272 131356 88324
rect 152464 88272 152516 88324
rect 411260 88272 411312 88324
rect 439964 88272 440016 88324
rect 131212 88204 131264 88256
rect 151268 88204 151320 88256
rect 423128 88204 423180 88256
rect 437480 88204 437532 88256
rect 132040 86980 132092 87032
rect 186320 86980 186372 87032
rect 131120 86912 131172 86964
rect 187148 86912 187200 86964
rect 411260 86912 411312 86964
rect 439872 86912 439924 86964
rect 131212 86844 131264 86896
rect 148416 86844 148468 86896
rect 425888 86844 425940 86896
rect 437480 86844 437532 86896
rect 133420 85552 133472 85604
rect 186320 85552 186372 85604
rect 540428 85552 540480 85604
rect 580172 85552 580224 85604
rect 132224 85484 132276 85536
rect 152556 85484 152608 85536
rect 423036 85484 423088 85536
rect 437480 85484 437532 85536
rect 131120 85416 131172 85468
rect 148508 85416 148560 85468
rect 132224 84804 132276 84856
rect 142896 84804 142948 84856
rect 131212 84124 131264 84176
rect 152648 84124 152700 84176
rect 131120 84056 131172 84108
rect 148600 84056 148652 84108
rect 142896 82900 142948 82952
rect 186320 82900 186372 82952
rect 135996 82832 136048 82884
rect 186412 82832 186464 82884
rect 411260 82832 411312 82884
rect 438216 82832 438268 82884
rect 131580 82764 131632 82816
rect 187240 82764 187292 82816
rect 417516 82764 417568 82816
rect 437480 82764 437532 82816
rect 131212 82696 131264 82748
rect 152740 82696 152792 82748
rect 132224 81336 132276 81388
rect 148692 81336 148744 81388
rect 422944 81336 422996 81388
rect 437480 81336 437532 81388
rect 131212 81268 131264 81320
rect 142988 81268 143040 81320
rect 411260 80112 411312 80164
rect 413560 80112 413612 80164
rect 136088 80044 136140 80096
rect 186320 80044 186372 80096
rect 131212 79976 131264 80028
rect 151360 79976 151412 80028
rect 417608 79976 417660 80028
rect 437480 79976 437532 80028
rect 131120 79908 131172 79960
rect 147220 79908 147272 79960
rect 131212 79840 131264 79892
rect 143080 79840 143132 79892
rect 138756 78684 138808 78736
rect 186320 78684 186372 78736
rect 131212 78616 131264 78668
rect 151084 78616 151136 78668
rect 421656 78616 421708 78668
rect 437480 78616 437532 78668
rect 131120 78548 131172 78600
rect 145564 78548 145616 78600
rect 411260 78276 411312 78328
rect 413652 78276 413704 78328
rect 131304 77936 131356 77988
rect 187332 77936 187384 77988
rect 131212 77188 131264 77240
rect 149704 77188 149756 77240
rect 411260 77188 411312 77240
rect 438124 77188 438176 77240
rect 131120 77120 131172 77172
rect 145748 77120 145800 77172
rect 138848 75964 138900 76016
rect 186320 75964 186372 76016
rect 134800 75896 134852 75948
rect 186412 75896 186464 75948
rect 131212 75828 131264 75880
rect 142804 75828 142856 75880
rect 419172 75828 419224 75880
rect 437480 75828 437532 75880
rect 131120 75760 131172 75812
rect 135904 75760 135956 75812
rect 159364 75216 159416 75268
rect 187516 75216 187568 75268
rect 132500 75148 132552 75200
rect 186964 75148 187016 75200
rect 131212 74468 131264 74520
rect 145656 74468 145708 74520
rect 411260 74468 411312 74520
rect 435548 74468 435600 74520
rect 131120 74400 131172 74452
rect 141792 74400 141844 74452
rect 421564 74400 421616 74452
rect 437480 74400 437532 74452
rect 132316 73176 132368 73228
rect 186320 73176 186372 73228
rect 131120 73108 131172 73160
rect 133696 73108 133748 73160
rect 429936 73108 429988 73160
rect 437480 73108 437532 73160
rect 131212 72972 131264 73024
rect 149796 72972 149848 73024
rect 411260 72768 411312 72820
rect 413468 72768 413520 72820
rect 181536 71748 181588 71800
rect 186320 71748 186372 71800
rect 131212 71680 131264 71732
rect 146944 71680 146996 71732
rect 417700 71680 417752 71732
rect 437480 71680 437532 71732
rect 131120 71612 131172 71664
rect 134524 71612 134576 71664
rect 133512 70388 133564 70440
rect 186320 70388 186372 70440
rect 131120 70320 131172 70372
rect 147036 70320 147088 70372
rect 426072 70320 426124 70372
rect 437480 70320 437532 70372
rect 131212 70252 131264 70304
rect 141424 70252 141476 70304
rect 146944 69096 146996 69148
rect 186412 69096 186464 69148
rect 134524 69028 134576 69080
rect 186320 69028 186372 69080
rect 131120 68960 131172 69012
rect 147128 68960 147180 69012
rect 131304 68892 131356 68944
rect 141516 68892 141568 68944
rect 131212 68824 131264 68876
rect 140044 68824 140096 68876
rect 181628 67600 181680 67652
rect 186320 67600 186372 67652
rect 411352 67600 411404 67652
rect 439872 67600 439924 67652
rect 131120 67532 131172 67584
rect 140136 67532 140188 67584
rect 411260 67532 411312 67584
rect 439780 67532 439832 67584
rect 425980 67464 426032 67516
rect 437480 67464 437532 67516
rect 131212 67328 131264 67380
rect 134616 67328 134668 67380
rect 144276 66240 144328 66292
rect 186320 66240 186372 66292
rect 131120 66172 131172 66224
rect 144184 66172 144236 66224
rect 431316 66172 431368 66224
rect 437480 66172 437532 66224
rect 131212 66104 131264 66156
rect 134708 66104 134760 66156
rect 411260 65016 411312 65068
rect 413468 65016 413520 65068
rect 134616 64880 134668 64932
rect 186320 64880 186372 64932
rect 131212 64812 131264 64864
rect 141608 64812 141660 64864
rect 424508 64812 424560 64864
rect 437480 64812 437532 64864
rect 131120 64744 131172 64796
rect 140228 64744 140280 64796
rect 181812 63520 181864 63572
rect 186320 63520 186372 63572
rect 132224 63452 132276 63504
rect 140320 63452 140372 63504
rect 411260 63452 411312 63504
rect 420276 63452 420328 63504
rect 142804 62092 142856 62144
rect 186320 62092 186372 62144
rect 131212 62024 131264 62076
rect 133236 62024 133288 62076
rect 424600 62024 424652 62076
rect 437480 62024 437532 62076
rect 132132 61956 132184 62008
rect 159364 61956 159416 62008
rect 131120 61888 131172 61940
rect 181444 61888 181496 61940
rect 181720 60800 181772 60852
rect 186320 60800 186372 60852
rect 134708 60732 134760 60784
rect 186412 60732 186464 60784
rect 411260 60732 411312 60784
rect 439780 60732 439832 60784
rect 131672 60664 131724 60716
rect 138664 60664 138716 60716
rect 411352 60664 411404 60716
rect 420184 60664 420236 60716
rect 540336 60664 540388 60716
rect 580172 60664 580224 60716
rect 132224 60596 132276 60648
rect 133328 60596 133380 60648
rect 141424 59372 141476 59424
rect 186320 59372 186372 59424
rect 131304 59304 131356 59356
rect 133420 59304 133472 59356
rect 432696 59304 432748 59356
rect 437480 59304 437532 59356
rect 133236 57944 133288 57996
rect 186320 57944 186372 57996
rect 131212 57876 131264 57928
rect 187056 57876 187108 57928
rect 416044 57876 416096 57928
rect 437480 57876 437532 57928
rect 131120 57808 131172 57860
rect 142896 57808 142948 57860
rect 411260 57808 411312 57860
rect 419080 57808 419132 57860
rect 131212 57740 131264 57792
rect 135996 57740 136048 57792
rect 132224 56516 132276 56568
rect 187148 56516 187200 56568
rect 435456 56516 435508 56568
rect 437756 56516 437808 56568
rect 131212 56448 131264 56500
rect 136088 56448 136140 56500
rect 132500 55836 132552 55888
rect 187424 55836 187476 55888
rect 140044 55224 140096 55276
rect 186320 55224 186372 55276
rect 411260 55224 411312 55276
rect 439964 55224 440016 55276
rect 131212 55156 131264 55208
rect 138756 55156 138808 55208
rect 416136 55156 416188 55208
rect 437480 55156 437532 55208
rect 131304 55088 131356 55140
rect 134800 55088 134852 55140
rect 133328 53796 133380 53848
rect 186320 53796 186372 53848
rect 131120 53728 131172 53780
rect 187240 53728 187292 53780
rect 424692 53728 424744 53780
rect 437480 53728 437532 53780
rect 131212 53660 131264 53712
rect 138848 53660 138900 53712
rect 131856 52436 131908 52488
rect 186320 52436 186372 52488
rect 131212 52368 131264 52420
rect 181536 52368 181588 52420
rect 133420 51076 133472 51128
rect 186320 51076 186372 51128
rect 131120 51008 131172 51060
rect 146944 51008 146996 51060
rect 131212 50940 131264 50992
rect 133512 50940 133564 50992
rect 411260 50940 411312 50992
rect 414756 50940 414808 50992
rect 131304 50872 131356 50924
rect 134524 50872 134576 50924
rect 131212 49648 131264 49700
rect 181628 49648 181680 49700
rect 423220 49648 423272 49700
rect 437480 49648 437532 49700
rect 131120 49580 131172 49632
rect 144276 49580 144328 49632
rect 132040 48288 132092 48340
rect 186320 48288 186372 48340
rect 131212 48220 131264 48272
rect 181812 48220 181864 48272
rect 411996 48220 412048 48272
rect 437480 48220 437532 48272
rect 131948 48016 132000 48068
rect 134616 48016 134668 48068
rect 411260 48016 411312 48068
rect 414848 48016 414900 48068
rect 132500 46928 132552 46980
rect 186320 46928 186372 46980
rect 131212 46860 131264 46912
rect 142804 46860 142856 46912
rect 421840 46860 421892 46912
rect 437480 46860 437532 46912
rect 131120 46792 131172 46844
rect 134708 46792 134760 46844
rect 411260 45568 411312 45620
rect 440056 45568 440108 45620
rect 540336 45568 540388 45620
rect 580172 45568 580224 45620
rect 131304 45500 131356 45552
rect 133236 45500 133288 45552
rect 421748 45500 421800 45552
rect 437480 45500 437532 45552
rect 131120 45432 131172 45484
rect 141424 45432 141476 45484
rect 131212 45364 131264 45416
rect 181720 45364 181772 45416
rect 182088 44140 182140 44192
rect 186320 44140 186372 44192
rect 131212 44072 131264 44124
rect 186964 44072 187016 44124
rect 131120 44004 131172 44056
rect 140044 44004 140096 44056
rect 131304 42780 131356 42832
rect 186320 42780 186372 42832
rect 131120 42712 131172 42764
rect 187056 42712 187108 42764
rect 411904 42712 411956 42764
rect 437480 42712 437532 42764
rect 131212 42644 131264 42696
rect 133328 42644 133380 42696
rect 411260 42508 411312 42560
rect 414664 42508 414716 42560
rect 131120 41352 131172 41404
rect 187148 41352 187200 41404
rect 411260 41352 411312 41404
rect 439688 41352 439740 41404
rect 131212 41284 131264 41336
rect 133420 41284 133472 41336
rect 417792 41284 417844 41336
rect 437480 41284 437532 41336
rect 413376 39992 413428 40044
rect 437480 39992 437532 40044
rect 131488 39312 131540 39364
rect 182088 39312 182140 39364
rect 131856 38632 131908 38684
rect 186320 38632 186372 38684
rect 131212 38564 131264 38616
rect 187424 38564 187476 38616
rect 411260 38564 411312 38616
rect 413284 38564 413336 38616
rect 418988 38564 419040 38616
rect 437480 38564 437532 38616
rect 131120 38496 131172 38548
rect 187240 38496 187292 38548
rect 132132 37272 132184 37324
rect 186320 37272 186372 37324
rect 131212 37204 131264 37256
rect 186412 37204 186464 37256
rect 411260 37204 411312 37256
rect 439596 37204 439648 37256
rect 132224 35912 132276 35964
rect 186320 35912 186372 35964
rect 131212 35844 131264 35896
rect 186964 35844 187016 35896
rect 417424 35844 417476 35896
rect 437480 35844 437532 35896
rect 131120 35776 131172 35828
rect 187056 35776 187108 35828
rect 411260 35776 411312 35828
rect 418804 35776 418856 35828
rect 414940 34416 414992 34468
rect 437480 34416 437532 34468
rect 131120 33124 131172 33176
rect 186320 33124 186372 33176
rect 131212 33056 131264 33108
rect 186412 33056 186464 33108
rect 412088 33056 412140 33108
rect 437480 33056 437532 33108
rect 411260 32988 411312 33040
rect 418896 32988 418948 33040
rect 131212 31832 131264 31884
rect 186412 31832 186464 31884
rect 131304 31764 131356 31816
rect 186320 31764 186372 31816
rect 411812 31696 411864 31748
rect 542728 31696 542780 31748
rect 412272 31628 412324 31680
rect 542544 31628 542596 31680
rect 412364 31560 412416 31612
rect 542636 31560 542688 31612
rect 412180 31492 412232 31544
rect 437480 31492 437532 31544
rect 131120 31016 131172 31068
rect 186320 31016 186372 31068
rect 439780 30268 439832 30320
rect 542452 30268 542504 30320
rect 439872 30200 439924 30252
rect 542360 30200 542412 30252
rect 131764 29248 131816 29300
rect 283012 29248 283064 29300
rect 440056 29248 440108 29300
rect 484584 29248 484636 29300
rect 130384 29180 130436 29232
rect 316224 29180 316276 29232
rect 438216 29180 438268 29232
rect 524604 29180 524656 29232
rect 206284 29112 206336 29164
rect 410524 29112 410576 29164
rect 435364 29112 435416 29164
rect 534632 29112 534684 29164
rect 130476 29044 130528 29096
rect 371240 29044 371292 29096
rect 413560 29044 413612 29096
rect 514760 29044 514812 29096
rect 205640 28976 205692 29028
rect 206284 28976 206336 29028
rect 217784 28976 217836 29028
rect 540336 28976 540388 29028
rect 79968 28908 80020 28960
rect 464620 28908 464672 28960
rect 195244 28840 195296 28892
rect 439504 28840 439556 28892
rect 445300 28840 445352 28892
rect 540428 28840 540480 28892
rect 188528 28772 188580 28824
rect 404452 28772 404504 28824
rect 413468 28772 413520 28824
rect 504640 28772 504692 28824
rect 188436 28704 188488 28756
rect 393412 28704 393464 28756
rect 455236 28704 455288 28756
rect 541624 28704 541676 28756
rect 166264 28636 166316 28688
rect 360200 28636 360252 28688
rect 411260 28636 411312 28688
rect 474740 28636 474792 28688
rect 190000 28568 190052 28620
rect 382280 28568 382332 28620
rect 439964 28568 440016 28620
rect 494612 28568 494664 28620
rect 164884 28500 164936 28552
rect 349160 28500 349212 28552
rect 188344 28432 188396 28484
rect 338120 28432 338172 28484
rect 189908 28364 189960 28416
rect 327080 28364 327132 28416
rect 133144 28296 133196 28348
rect 239036 28296 239088 28348
rect 190092 28228 190144 28280
rect 294052 28228 294104 28280
rect 189724 28160 189776 28212
rect 271972 28160 272024 28212
rect 189816 28092 189868 28144
rect 261116 28092 261168 28144
rect 190184 28024 190236 28076
rect 250076 28024 250128 28076
rect 540244 20612 540296 20664
rect 579988 20612 580040 20664
rect 227720 6808 227772 6860
rect 580172 6808 580224 6860
rect 2688 4088 2740 4140
rect 205640 4088 205692 4140
rect 1308 4020 1360 4072
rect 195244 4020 195296 4072
rect 1676 3680 1728 3732
rect 2688 3680 2740 3732
rect 572 3612 624 3664
rect 1308 3612 1360 3664
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 48226 334248 48282 334257
rect 48226 334183 48282 334192
rect 47766 333024 47822 333033
rect 47766 332959 47822 332968
rect 47674 330168 47730 330177
rect 47674 330103 47730 330112
rect 47688 279478 47716 330103
rect 47780 287706 47808 332959
rect 47858 331120 47914 331129
rect 47858 331055 47914 331064
rect 47768 287700 47820 287706
rect 47768 287642 47820 287648
rect 47872 282198 47900 331055
rect 48134 325816 48190 325825
rect 48134 325751 48190 325760
rect 48042 307320 48098 307329
rect 48042 307255 48098 307264
rect 47860 282192 47912 282198
rect 47860 282134 47912 282140
rect 47676 279472 47728 279478
rect 47676 279414 47728 279420
rect 1308 131232 1360 131238
rect 1308 131174 1360 131180
rect 1320 4078 1348 131174
rect 2688 131164 2740 131170
rect 2688 131106 2740 131112
rect 2700 4146 2728 131106
rect 48056 130558 48084 307255
rect 48148 131782 48176 325751
rect 48136 131776 48188 131782
rect 48136 131718 48188 131724
rect 48044 130552 48096 130558
rect 48044 130494 48096 130500
rect 48240 130422 48268 334183
rect 209686 334112 209742 334121
rect 209686 334047 209742 334056
rect 208306 332888 208362 332897
rect 208306 332823 208362 332832
rect 208214 331120 208270 331129
rect 208214 331055 208270 331064
rect 49606 328490 49662 328499
rect 49606 328425 49662 328434
rect 49514 327538 49570 327547
rect 49514 327473 49570 327482
rect 49422 305642 49478 305651
rect 49422 305577 49478 305586
rect 49436 291854 49464 305577
rect 49424 291848 49476 291854
rect 49424 291790 49476 291796
rect 49528 279546 49556 327473
rect 49516 279540 49568 279546
rect 49516 279482 49568 279488
rect 49620 233238 49648 328425
rect 208122 327448 208178 327457
rect 208122 327383 208178 327392
rect 207018 325816 207074 325825
rect 207018 325751 207074 325760
rect 207032 325718 207060 325751
rect 204260 325712 204312 325718
rect 204260 325654 204312 325660
rect 207020 325712 207072 325718
rect 207020 325654 207072 325660
rect 193220 306400 193272 306406
rect 193220 306342 193272 306348
rect 190460 305040 190512 305046
rect 190460 304982 190512 304988
rect 55862 299568 55918 299577
rect 55862 299503 55918 299512
rect 67822 299568 67878 299577
rect 67822 299503 67878 299512
rect 55876 298178 55904 299503
rect 67836 298314 67864 299503
rect 67824 298308 67876 298314
rect 67824 298250 67876 298256
rect 69296 298240 69348 298246
rect 69296 298182 69348 298188
rect 55220 298172 55272 298178
rect 55220 298114 55272 298120
rect 55864 298172 55916 298178
rect 55864 298114 55916 298120
rect 49608 233232 49660 233238
rect 49608 233174 49660 233180
rect 55128 131232 55180 131238
rect 55232 131186 55260 298114
rect 69308 298081 69336 298182
rect 65798 298072 65854 298081
rect 65798 298007 65854 298016
rect 67546 298072 67602 298081
rect 67546 298007 67602 298016
rect 69294 298072 69350 298081
rect 69294 298007 69350 298016
rect 70214 298072 70270 298081
rect 70214 298007 70270 298016
rect 71686 298072 71742 298081
rect 71686 298007 71742 298016
rect 73066 298072 73122 298081
rect 73066 298007 73122 298016
rect 74446 298072 74502 298081
rect 74446 298007 74502 298016
rect 75550 298072 75606 298081
rect 75550 298007 75606 298016
rect 76838 298072 76894 298081
rect 76838 298007 76840 298016
rect 65812 296750 65840 298007
rect 65800 296744 65852 296750
rect 65800 296686 65852 296692
rect 67560 252550 67588 298007
rect 70228 297294 70256 298007
rect 70216 297288 70268 297294
rect 70216 297230 70268 297236
rect 67548 252544 67600 252550
rect 67548 252486 67600 252492
rect 71700 230450 71728 298007
rect 73080 231810 73108 298007
rect 74460 260370 74488 298007
rect 75564 297362 75592 298007
rect 76892 298007 76894 298016
rect 77114 298072 77170 298081
rect 77114 298007 77170 298016
rect 78494 298072 78550 298081
rect 79874 298072 79930 298081
rect 78494 298007 78550 298016
rect 79324 298036 79376 298042
rect 76840 297978 76892 297984
rect 75552 297356 75604 297362
rect 75552 297298 75604 297304
rect 74448 260364 74500 260370
rect 74448 260306 74500 260312
rect 77128 251870 77156 298007
rect 77116 251864 77168 251870
rect 77116 251806 77168 251812
rect 78508 250510 78536 298007
rect 79874 298007 79930 298016
rect 81254 298072 81310 298081
rect 81254 298007 81310 298016
rect 82634 298072 82690 298081
rect 82634 298007 82690 298016
rect 84014 298072 84070 298081
rect 84014 298007 84070 298016
rect 85486 298072 85542 298081
rect 85486 298007 85542 298016
rect 86682 298072 86738 298081
rect 86682 298007 86738 298016
rect 88154 298072 88210 298081
rect 88154 298007 88210 298016
rect 89166 298072 89222 298081
rect 89166 298007 89222 298016
rect 89534 298072 89590 298081
rect 89534 298007 89590 298016
rect 91006 298072 91062 298081
rect 91006 298007 91062 298016
rect 92294 298072 92350 298081
rect 92294 298007 92350 298016
rect 93674 298072 93730 298081
rect 93674 298007 93730 298016
rect 95054 298072 95110 298081
rect 95054 298007 95110 298016
rect 96434 298072 96490 298081
rect 96434 298007 96490 298016
rect 97078 298072 97134 298081
rect 97078 298007 97134 298016
rect 97906 298072 97962 298081
rect 97906 298007 97962 298016
rect 100666 298072 100722 298081
rect 100666 298007 100722 298016
rect 101862 298072 101918 298081
rect 101862 298007 101918 298016
rect 102966 298072 103022 298081
rect 102966 298007 103022 298016
rect 103334 298072 103390 298081
rect 103334 298007 103390 298016
rect 104254 298072 104310 298081
rect 104254 298007 104310 298016
rect 104714 298072 104770 298081
rect 104714 298007 104770 298016
rect 105542 298072 105598 298081
rect 105542 298007 105598 298016
rect 106094 298072 106150 298081
rect 106094 298007 106150 298016
rect 106646 298072 106702 298081
rect 106646 298007 106702 298016
rect 107474 298072 107530 298081
rect 107474 298007 107530 298016
rect 107750 298072 107806 298081
rect 107750 298007 107806 298016
rect 108854 298072 108910 298081
rect 108854 298007 108910 298016
rect 110326 298072 110382 298081
rect 110326 298007 110382 298016
rect 111614 298072 111670 298081
rect 111614 298007 111670 298016
rect 112994 298072 113050 298081
rect 112994 298007 113050 298016
rect 114466 298072 114522 298081
rect 114466 298007 114522 298016
rect 115846 298072 115902 298081
rect 115846 298007 115902 298016
rect 117226 298072 117282 298081
rect 117226 298007 117282 298016
rect 79324 297978 79376 297984
rect 78586 297936 78642 297945
rect 78586 297871 78642 297880
rect 78496 250504 78548 250510
rect 78496 250446 78548 250452
rect 73068 231804 73120 231810
rect 73068 231746 73120 231752
rect 71688 230444 71740 230450
rect 71688 230386 71740 230392
rect 55180 131180 55260 131186
rect 55128 131174 55260 131180
rect 55140 131158 55260 131174
rect 48228 130416 48280 130422
rect 48228 130358 48280 130364
rect 55140 129962 55168 131158
rect 78600 130490 78628 297871
rect 79336 251938 79364 297978
rect 79888 260302 79916 298007
rect 79966 297936 80022 297945
rect 79966 297871 80022 297880
rect 79876 260296 79928 260302
rect 79876 260238 79928 260244
rect 79324 251932 79376 251938
rect 79324 251874 79376 251880
rect 79980 191146 80008 297871
rect 81268 262886 81296 298007
rect 81346 297936 81402 297945
rect 81346 297871 81402 297880
rect 81256 262880 81308 262886
rect 81256 262822 81308 262828
rect 81360 257378 81388 297871
rect 81348 257372 81400 257378
rect 81348 257314 81400 257320
rect 82648 254590 82676 298007
rect 82726 297936 82782 297945
rect 82726 297871 82782 297880
rect 82636 254584 82688 254590
rect 82636 254526 82688 254532
rect 82740 250578 82768 297871
rect 84028 256018 84056 298007
rect 84106 297936 84162 297945
rect 84106 297871 84162 297880
rect 85394 297936 85450 297945
rect 85394 297871 85450 297880
rect 84016 256012 84068 256018
rect 84016 255954 84068 255960
rect 82728 250572 82780 250578
rect 82728 250514 82780 250520
rect 84120 237386 84148 297871
rect 85302 297120 85358 297129
rect 85302 297055 85358 297064
rect 85316 279614 85344 297055
rect 85304 279608 85356 279614
rect 85304 279550 85356 279556
rect 85408 258738 85436 297871
rect 85396 258732 85448 258738
rect 85396 258674 85448 258680
rect 85500 246362 85528 298007
rect 86696 261526 86724 298007
rect 86774 297936 86830 297945
rect 86774 297871 86830 297880
rect 86684 261520 86736 261526
rect 86684 261462 86736 261468
rect 85488 246356 85540 246362
rect 85488 246298 85540 246304
rect 84108 237380 84160 237386
rect 84108 237322 84160 237328
rect 86788 234598 86816 297871
rect 86866 297800 86922 297809
rect 86866 297735 86922 297744
rect 86776 234592 86828 234598
rect 86776 234534 86828 234540
rect 86880 233170 86908 297735
rect 88168 261662 88196 298007
rect 88246 297936 88302 297945
rect 88246 297871 88302 297880
rect 88156 261656 88208 261662
rect 88156 261598 88208 261604
rect 88260 241466 88288 297871
rect 89180 297430 89208 298007
rect 89168 297424 89220 297430
rect 89168 297366 89220 297372
rect 88248 241460 88300 241466
rect 88248 241402 88300 241408
rect 89548 235958 89576 298007
rect 90914 297936 90970 297945
rect 90914 297871 90970 297880
rect 90928 261594 90956 297871
rect 90916 261588 90968 261594
rect 90916 261530 90968 261536
rect 91020 254658 91048 298007
rect 92308 254726 92336 298007
rect 92386 297936 92442 297945
rect 92386 297871 92442 297880
rect 93582 297936 93638 297945
rect 93582 297871 93638 297880
rect 92296 254720 92348 254726
rect 92296 254662 92348 254668
rect 91008 254652 91060 254658
rect 91008 254594 91060 254600
rect 89536 235952 89588 235958
rect 89536 235894 89588 235900
rect 86868 233164 86920 233170
rect 86868 233106 86920 233112
rect 92400 191214 92428 297871
rect 93596 258806 93624 297871
rect 93584 258800 93636 258806
rect 93584 258742 93636 258748
rect 93688 191282 93716 298007
rect 93766 297800 93822 297809
rect 93766 297735 93822 297744
rect 93676 191276 93728 191282
rect 93676 191218 93728 191224
rect 92388 191208 92440 191214
rect 92388 191150 92440 191156
rect 79968 191140 80020 191146
rect 79968 191082 80020 191088
rect 93780 133346 93808 297735
rect 95068 247042 95096 298007
rect 95146 297936 95202 297945
rect 95146 297871 95202 297880
rect 95056 247036 95108 247042
rect 95056 246978 95108 246984
rect 95160 240106 95188 297871
rect 96448 262954 96476 298007
rect 96526 297936 96582 297945
rect 96526 297871 96582 297880
rect 96436 262948 96488 262954
rect 96436 262890 96488 262896
rect 95148 240100 95200 240106
rect 95148 240042 95200 240048
rect 96540 240038 96568 297871
rect 97092 297498 97120 298007
rect 97814 297936 97870 297945
rect 97814 297871 97870 297880
rect 97080 297492 97132 297498
rect 97080 297434 97132 297440
rect 97828 256086 97856 297871
rect 97816 256080 97868 256086
rect 97816 256022 97868 256028
rect 96528 240032 96580 240038
rect 96528 239974 96580 239980
rect 93768 133340 93820 133346
rect 93768 133282 93820 133288
rect 97920 131850 97948 298007
rect 100574 297936 100630 297945
rect 100574 297871 100630 297880
rect 100588 264246 100616 297871
rect 100576 264240 100628 264246
rect 100576 264182 100628 264188
rect 100680 242894 100708 298007
rect 101876 244254 101904 298007
rect 101954 297936 102010 297945
rect 101954 297871 102010 297880
rect 101968 250646 101996 297871
rect 102046 297800 102102 297809
rect 102046 297735 102102 297744
rect 102060 296818 102088 297735
rect 102980 296886 103008 298007
rect 102968 296880 103020 296886
rect 102968 296822 103020 296828
rect 102048 296812 102100 296818
rect 102048 296754 102100 296760
rect 101956 250640 102008 250646
rect 101956 250582 102008 250588
rect 103348 245614 103376 298007
rect 104268 296954 104296 298007
rect 104256 296948 104308 296954
rect 104256 296890 104308 296896
rect 104728 257446 104756 298007
rect 105556 297022 105584 298007
rect 105544 297016 105596 297022
rect 105544 296958 105596 296964
rect 104716 257440 104768 257446
rect 104716 257382 104768 257388
rect 106108 248402 106136 298007
rect 106660 297226 106688 298007
rect 106648 297220 106700 297226
rect 106648 297162 106700 297168
rect 106096 248396 106148 248402
rect 106096 248338 106148 248344
rect 107488 248334 107516 298007
rect 107764 297158 107792 298007
rect 107752 297152 107804 297158
rect 107752 297094 107804 297100
rect 108868 257514 108896 298007
rect 108856 257508 108908 257514
rect 108856 257450 108908 257456
rect 107476 248328 107528 248334
rect 107476 248270 107528 248276
rect 103336 245608 103388 245614
rect 103336 245550 103388 245556
rect 101864 244248 101916 244254
rect 101864 244190 101916 244196
rect 100668 242888 100720 242894
rect 100668 242830 100720 242836
rect 110340 131918 110368 298007
rect 111628 297090 111656 298007
rect 111616 297084 111668 297090
rect 111616 297026 111668 297032
rect 113008 260166 113036 298007
rect 113086 297936 113142 297945
rect 113086 297871 113142 297880
rect 112996 260160 113048 260166
rect 112996 260102 113048 260108
rect 113100 133210 113128 297871
rect 114480 249762 114508 298007
rect 115860 260234 115888 298007
rect 115848 260228 115900 260234
rect 115848 260170 115900 260176
rect 114468 249756 114520 249762
rect 114468 249698 114520 249704
rect 117240 133278 117268 298007
rect 130476 297492 130528 297498
rect 130476 297434 130528 297440
rect 130384 297424 130436 297430
rect 130384 297366 130436 297372
rect 117228 133272 117280 133278
rect 117228 133214 117280 133220
rect 113088 133204 113140 133210
rect 113088 133146 113140 133152
rect 110328 131912 110380 131918
rect 110328 131854 110380 131860
rect 97908 131844 97960 131850
rect 97908 131786 97960 131792
rect 104900 131164 104952 131170
rect 104900 131106 104952 131112
rect 78588 130484 78640 130490
rect 78588 130426 78640 130432
rect 54978 129934 55168 129962
rect 104912 129948 104940 131106
rect 79980 28966 80008 30056
rect 130396 29238 130424 297366
rect 130384 29232 130436 29238
rect 130384 29174 130436 29180
rect 130488 29102 130516 297434
rect 131764 297356 131816 297362
rect 131764 297298 131816 297304
rect 131120 129736 131172 129742
rect 131118 129704 131120 129713
rect 131172 129704 131174 129713
rect 131118 129639 131174 129648
rect 131304 129668 131356 129674
rect 131304 129610 131356 129616
rect 131212 129600 131264 129606
rect 131212 129542 131264 129548
rect 131224 129169 131252 129542
rect 131210 129160 131266 129169
rect 131210 129095 131266 129104
rect 131316 128625 131344 129610
rect 131302 128616 131358 128625
rect 131302 128551 131358 128560
rect 131120 126948 131172 126954
rect 131120 126890 131172 126896
rect 131132 126177 131160 126890
rect 131210 126848 131266 126857
rect 131210 126783 131212 126792
rect 131264 126783 131266 126792
rect 131212 126754 131264 126760
rect 131118 126168 131174 126177
rect 131118 126103 131174 126112
rect 131120 125588 131172 125594
rect 131120 125530 131172 125536
rect 131132 125089 131160 125530
rect 131212 125520 131264 125526
rect 131212 125462 131264 125468
rect 131118 125080 131174 125089
rect 131118 125015 131174 125024
rect 131224 124545 131252 125462
rect 131210 124536 131266 124545
rect 131210 124471 131266 124480
rect 131120 124092 131172 124098
rect 131120 124034 131172 124040
rect 131132 123321 131160 124034
rect 131118 123312 131174 123321
rect 131118 123247 131174 123256
rect 131212 122800 131264 122806
rect 131210 122768 131212 122777
rect 131264 122768 131266 122777
rect 131120 122732 131172 122738
rect 131210 122703 131266 122712
rect 131120 122674 131172 122680
rect 131132 121553 131160 122674
rect 131212 122664 131264 122670
rect 131212 122606 131264 122612
rect 131224 122097 131252 122606
rect 131210 122088 131266 122097
rect 131210 122023 131266 122032
rect 131118 121544 131174 121553
rect 131118 121479 131174 121488
rect 131212 121372 131264 121378
rect 131212 121314 131264 121320
rect 131224 121009 131252 121314
rect 131210 121000 131266 121009
rect 131210 120935 131266 120944
rect 131120 120012 131172 120018
rect 131120 119954 131172 119960
rect 131132 119241 131160 119954
rect 131118 119232 131174 119241
rect 131118 119167 131174 119176
rect 131210 118688 131266 118697
rect 131210 118623 131212 118632
rect 131264 118623 131266 118632
rect 131212 118594 131264 118600
rect 131120 118584 131172 118590
rect 131120 118526 131172 118532
rect 131132 118017 131160 118526
rect 131212 118516 131264 118522
rect 131212 118458 131264 118464
rect 131118 118008 131174 118017
rect 131118 117943 131174 117952
rect 131224 117473 131252 118458
rect 131210 117464 131266 117473
rect 131210 117399 131266 117408
rect 131212 117292 131264 117298
rect 131212 117234 131264 117240
rect 131120 117224 131172 117230
rect 131120 117166 131172 117172
rect 131132 116249 131160 117166
rect 131224 116929 131252 117234
rect 131210 116920 131266 116929
rect 131210 116855 131266 116864
rect 131118 116240 131174 116249
rect 131118 116175 131174 116184
rect 131212 115932 131264 115938
rect 131212 115874 131264 115880
rect 131224 115705 131252 115874
rect 131210 115696 131266 115705
rect 131210 115631 131266 115640
rect 131212 115524 131264 115530
rect 131212 115466 131264 115472
rect 131224 115161 131252 115466
rect 131210 115152 131266 115161
rect 131210 115087 131266 115096
rect 131304 114504 131356 114510
rect 131210 114472 131266 114481
rect 131304 114446 131356 114452
rect 131210 114407 131212 114416
rect 131264 114407 131266 114416
rect 131212 114378 131264 114384
rect 131120 114368 131172 114374
rect 131120 114310 131172 114316
rect 131132 113393 131160 114310
rect 131316 113937 131344 114446
rect 131302 113928 131358 113937
rect 131302 113863 131358 113872
rect 131118 113384 131174 113393
rect 131118 113319 131174 113328
rect 131212 113144 131264 113150
rect 131212 113086 131264 113092
rect 131120 113076 131172 113082
rect 131120 113018 131172 113024
rect 131132 112169 131160 113018
rect 131224 112849 131252 113086
rect 131210 112840 131266 112849
rect 131210 112775 131266 112784
rect 131118 112160 131174 112169
rect 131118 112095 131174 112104
rect 131212 111716 131264 111722
rect 131212 111658 131264 111664
rect 131224 111081 131252 111658
rect 131210 111072 131266 111081
rect 131210 111007 131266 111016
rect 131304 110424 131356 110430
rect 131210 110392 131266 110401
rect 131304 110366 131356 110372
rect 131210 110327 131212 110336
rect 131264 110327 131266 110336
rect 131212 110298 131264 110304
rect 131120 110288 131172 110294
rect 131120 110230 131172 110236
rect 131132 109857 131160 110230
rect 131118 109848 131174 109857
rect 131118 109783 131174 109792
rect 131316 109313 131344 110366
rect 131302 109304 131358 109313
rect 131302 109239 131358 109248
rect 131120 108996 131172 109002
rect 131120 108938 131172 108944
rect 131132 108089 131160 108938
rect 131212 108928 131264 108934
rect 131212 108870 131264 108876
rect 131224 108633 131252 108870
rect 131210 108624 131266 108633
rect 131210 108559 131266 108568
rect 131118 108080 131174 108089
rect 131118 108015 131174 108024
rect 131120 107636 131172 107642
rect 131120 107578 131172 107584
rect 131132 107001 131160 107578
rect 131304 107568 131356 107574
rect 131210 107536 131266 107545
rect 131304 107510 131356 107516
rect 131210 107471 131212 107480
rect 131264 107471 131266 107480
rect 131212 107442 131264 107448
rect 131118 106992 131174 107001
rect 131118 106927 131174 106936
rect 131316 106321 131344 107510
rect 131302 106312 131358 106321
rect 131120 106276 131172 106282
rect 131302 106247 131358 106256
rect 131120 106218 131172 106224
rect 131132 105777 131160 106218
rect 131212 106208 131264 106214
rect 131212 106150 131264 106156
rect 131118 105768 131174 105777
rect 131118 105703 131174 105712
rect 131224 105233 131252 106150
rect 131210 105224 131266 105233
rect 131210 105159 131266 105168
rect 131212 104848 131264 104854
rect 131212 104790 131264 104796
rect 131120 104780 131172 104786
rect 131120 104722 131172 104728
rect 131132 104009 131160 104722
rect 131224 104553 131252 104790
rect 131210 104544 131266 104553
rect 131210 104479 131266 104488
rect 131118 104000 131174 104009
rect 131118 103935 131174 103944
rect 131672 103488 131724 103494
rect 131210 103456 131266 103465
rect 131672 103430 131724 103436
rect 131210 103391 131212 103400
rect 131264 103391 131266 103400
rect 131212 103362 131264 103368
rect 131120 103352 131172 103358
rect 131120 103294 131172 103300
rect 131132 102241 131160 103294
rect 131684 102785 131712 103430
rect 131670 102776 131726 102785
rect 131670 102711 131726 102720
rect 131118 102232 131174 102241
rect 131118 102167 131174 102176
rect 131212 102128 131264 102134
rect 131212 102070 131264 102076
rect 131120 102060 131172 102066
rect 131120 102002 131172 102008
rect 131132 101153 131160 102002
rect 131224 101697 131252 102070
rect 131210 101688 131266 101697
rect 131210 101623 131266 101632
rect 131118 101144 131174 101153
rect 131118 101079 131174 101088
rect 131212 100700 131264 100706
rect 131212 100642 131264 100648
rect 131224 99929 131252 100642
rect 131488 100020 131540 100026
rect 131488 99962 131540 99968
rect 131210 99920 131266 99929
rect 131210 99855 131266 99864
rect 131210 99376 131266 99385
rect 131210 99311 131212 99320
rect 131264 99311 131266 99320
rect 131212 99282 131264 99288
rect 131120 99272 131172 99278
rect 131120 99214 131172 99220
rect 131132 98705 131160 99214
rect 131118 98696 131174 98705
rect 131118 98631 131174 98640
rect 131500 98161 131528 99962
rect 131486 98152 131542 98161
rect 131486 98087 131542 98096
rect 131120 97980 131172 97986
rect 131120 97922 131172 97928
rect 131132 97073 131160 97922
rect 131212 97912 131264 97918
rect 131212 97854 131264 97860
rect 131224 97617 131252 97854
rect 131210 97608 131266 97617
rect 131210 97543 131266 97552
rect 131118 97064 131174 97073
rect 131118 96999 131174 97008
rect 131120 96620 131172 96626
rect 131120 96562 131172 96568
rect 131132 95849 131160 96562
rect 131212 96484 131264 96490
rect 131212 96426 131264 96432
rect 131224 96393 131252 96426
rect 131210 96384 131266 96393
rect 131210 96319 131266 96328
rect 131118 95840 131174 95849
rect 131118 95775 131174 95784
rect 131212 95192 131264 95198
rect 131212 95134 131264 95140
rect 131120 95124 131172 95130
rect 131120 95066 131172 95072
rect 131132 94081 131160 95066
rect 131224 94625 131252 95134
rect 131210 94616 131266 94625
rect 131210 94551 131266 94560
rect 131118 94072 131174 94081
rect 131118 94007 131174 94016
rect 131212 93832 131264 93838
rect 131212 93774 131264 93780
rect 131120 93764 131172 93770
rect 131120 93706 131172 93712
rect 131132 92857 131160 93706
rect 131224 93537 131252 93774
rect 131210 93528 131266 93537
rect 131210 93463 131266 93472
rect 131118 92848 131174 92857
rect 131118 92783 131174 92792
rect 131304 92472 131356 92478
rect 131304 92414 131356 92420
rect 131120 92404 131172 92410
rect 131120 92346 131172 92352
rect 131132 91769 131160 92346
rect 131212 92336 131264 92342
rect 131210 92304 131212 92313
rect 131264 92304 131266 92313
rect 131210 92239 131266 92248
rect 131118 91760 131174 91769
rect 131118 91695 131174 91704
rect 131316 91225 131344 92414
rect 131302 91216 131358 91225
rect 131302 91151 131358 91160
rect 131212 91044 131264 91050
rect 131212 90986 131264 90992
rect 131120 90976 131172 90982
rect 131120 90918 131172 90924
rect 131132 90001 131160 90918
rect 131224 90545 131252 90986
rect 131210 90536 131266 90545
rect 131210 90471 131266 90480
rect 131118 89992 131174 90001
rect 131118 89927 131174 89936
rect 131304 89684 131356 89690
rect 131304 89626 131356 89632
rect 131120 89004 131172 89010
rect 131120 88946 131172 88952
rect 131132 87689 131160 88946
rect 131316 88777 131344 89626
rect 131302 88768 131358 88777
rect 131302 88703 131358 88712
rect 131304 88324 131356 88330
rect 131304 88266 131356 88272
rect 131212 88256 131264 88262
rect 131210 88224 131212 88233
rect 131264 88224 131266 88233
rect 131210 88159 131266 88168
rect 131118 87680 131174 87689
rect 131118 87615 131174 87624
rect 131316 87009 131344 88266
rect 131302 87000 131358 87009
rect 131120 86964 131172 86970
rect 131302 86935 131358 86944
rect 131120 86906 131172 86912
rect 131132 85921 131160 86906
rect 131212 86896 131264 86902
rect 131212 86838 131264 86844
rect 131224 86465 131252 86838
rect 131210 86456 131266 86465
rect 131210 86391 131266 86400
rect 131118 85912 131174 85921
rect 131118 85847 131174 85856
rect 131120 85468 131172 85474
rect 131120 85410 131172 85416
rect 131132 84697 131160 85410
rect 131118 84688 131174 84697
rect 131118 84623 131174 84632
rect 131212 84176 131264 84182
rect 131212 84118 131264 84124
rect 131120 84108 131172 84114
rect 131120 84050 131172 84056
rect 131132 82929 131160 84050
rect 131224 83609 131252 84118
rect 131210 83600 131266 83609
rect 131210 83535 131266 83544
rect 131118 82920 131174 82929
rect 131118 82855 131174 82864
rect 131580 82816 131632 82822
rect 131580 82758 131632 82764
rect 131212 82748 131264 82754
rect 131212 82690 131264 82696
rect 131224 81841 131252 82690
rect 131592 82385 131620 82758
rect 131578 82376 131634 82385
rect 131578 82311 131634 82320
rect 131210 81832 131266 81841
rect 131210 81767 131266 81776
rect 131212 81320 131264 81326
rect 131212 81262 131264 81268
rect 131224 80617 131252 81262
rect 131210 80608 131266 80617
rect 131210 80543 131266 80552
rect 131210 80064 131266 80073
rect 131210 79999 131212 80008
rect 131264 79999 131266 80008
rect 131212 79970 131264 79976
rect 131120 79960 131172 79966
rect 131120 79902 131172 79908
rect 131132 79529 131160 79902
rect 131212 79892 131264 79898
rect 131212 79834 131264 79840
rect 131118 79520 131174 79529
rect 131118 79455 131174 79464
rect 131224 78849 131252 79834
rect 131210 78840 131266 78849
rect 131210 78775 131266 78784
rect 131212 78668 131264 78674
rect 131212 78610 131264 78616
rect 131120 78600 131172 78606
rect 131120 78542 131172 78548
rect 131132 77761 131160 78542
rect 131224 78305 131252 78610
rect 131210 78296 131266 78305
rect 131210 78231 131266 78240
rect 131304 77988 131356 77994
rect 131304 77930 131356 77936
rect 131118 77752 131174 77761
rect 131118 77687 131174 77696
rect 131212 77240 131264 77246
rect 131212 77182 131264 77188
rect 131120 77172 131172 77178
rect 131120 77114 131172 77120
rect 131132 75993 131160 77114
rect 131224 76537 131252 77182
rect 131316 77081 131344 77930
rect 131302 77072 131358 77081
rect 131302 77007 131358 77016
rect 131210 76528 131266 76537
rect 131210 76463 131266 76472
rect 131118 75984 131174 75993
rect 131118 75919 131174 75928
rect 131212 75880 131264 75886
rect 131212 75822 131264 75828
rect 131120 75812 131172 75818
rect 131120 75754 131172 75760
rect 131132 74769 131160 75754
rect 131224 75313 131252 75822
rect 131210 75304 131266 75313
rect 131210 75239 131266 75248
rect 131118 74760 131174 74769
rect 131118 74695 131174 74704
rect 131212 74520 131264 74526
rect 131212 74462 131264 74468
rect 131120 74452 131172 74458
rect 131120 74394 131172 74400
rect 131132 73681 131160 74394
rect 131224 74225 131252 74462
rect 131210 74216 131266 74225
rect 131210 74151 131266 74160
rect 131118 73672 131174 73681
rect 131118 73607 131174 73616
rect 131120 73160 131172 73166
rect 131120 73102 131172 73108
rect 131132 72457 131160 73102
rect 131212 73024 131264 73030
rect 131210 72992 131212 73001
rect 131264 72992 131266 73001
rect 131210 72927 131266 72936
rect 131118 72448 131174 72457
rect 131118 72383 131174 72392
rect 131212 71732 131264 71738
rect 131212 71674 131264 71680
rect 131120 71664 131172 71670
rect 131120 71606 131172 71612
rect 131132 70689 131160 71606
rect 131224 71233 131252 71674
rect 131210 71224 131266 71233
rect 131210 71159 131266 71168
rect 131118 70680 131174 70689
rect 131118 70615 131174 70624
rect 131120 70372 131172 70378
rect 131120 70314 131172 70320
rect 131132 69465 131160 70314
rect 131212 70304 131264 70310
rect 131212 70246 131264 70252
rect 131224 70145 131252 70246
rect 131210 70136 131266 70145
rect 131210 70071 131266 70080
rect 131118 69456 131174 69465
rect 131118 69391 131174 69400
rect 131120 69012 131172 69018
rect 131120 68954 131172 68960
rect 131132 68921 131160 68954
rect 131304 68944 131356 68950
rect 131118 68912 131174 68921
rect 131304 68886 131356 68892
rect 131118 68847 131174 68856
rect 131212 68876 131264 68882
rect 131212 68818 131264 68824
rect 131224 68377 131252 68818
rect 131210 68368 131266 68377
rect 131210 68303 131266 68312
rect 131316 67833 131344 68886
rect 131302 67824 131358 67833
rect 131302 67759 131358 67768
rect 131120 67584 131172 67590
rect 131120 67526 131172 67532
rect 131132 66609 131160 67526
rect 131212 67380 131264 67386
rect 131212 67322 131264 67328
rect 131224 67153 131252 67322
rect 131210 67144 131266 67153
rect 131210 67079 131266 67088
rect 131118 66600 131174 66609
rect 131118 66535 131174 66544
rect 131120 66224 131172 66230
rect 131120 66166 131172 66172
rect 131132 65385 131160 66166
rect 131212 66156 131264 66162
rect 131212 66098 131264 66104
rect 131224 66065 131252 66098
rect 131210 66056 131266 66065
rect 131210 65991 131266 66000
rect 131118 65376 131174 65385
rect 131118 65311 131174 65320
rect 131212 64864 131264 64870
rect 131210 64832 131212 64841
rect 131264 64832 131266 64841
rect 131120 64796 131172 64802
rect 131210 64767 131266 64776
rect 131120 64738 131172 64744
rect 131132 63753 131160 64738
rect 131118 63744 131174 63753
rect 131118 63679 131174 63688
rect 131212 62076 131264 62082
rect 131212 62018 131264 62024
rect 131224 61985 131252 62018
rect 131210 61976 131266 61985
rect 131120 61940 131172 61946
rect 131210 61911 131266 61920
rect 131120 61882 131172 61888
rect 131132 60761 131160 61882
rect 131118 60752 131174 60761
rect 131118 60687 131174 60696
rect 131672 60716 131724 60722
rect 131672 60658 131724 60664
rect 131684 59537 131712 60658
rect 131670 59528 131726 59537
rect 131670 59463 131726 59472
rect 131304 59356 131356 59362
rect 131304 59298 131356 59304
rect 131316 58449 131344 59298
rect 131302 58440 131358 58449
rect 131302 58375 131358 58384
rect 131212 57928 131264 57934
rect 131210 57896 131212 57905
rect 131264 57896 131266 57905
rect 131120 57860 131172 57866
rect 131210 57831 131266 57840
rect 131120 57802 131172 57808
rect 131132 56681 131160 57802
rect 131212 57792 131264 57798
rect 131212 57734 131264 57740
rect 131224 57225 131252 57734
rect 131210 57216 131266 57225
rect 131210 57151 131266 57160
rect 131118 56672 131174 56681
rect 131118 56607 131174 56616
rect 131212 56500 131264 56506
rect 131212 56442 131264 56448
rect 131224 55457 131252 56442
rect 131210 55448 131266 55457
rect 131210 55383 131266 55392
rect 131212 55208 131264 55214
rect 131212 55150 131264 55156
rect 131224 54913 131252 55150
rect 131304 55140 131356 55146
rect 131304 55082 131356 55088
rect 131210 54904 131266 54913
rect 131210 54839 131266 54848
rect 131120 53780 131172 53786
rect 131120 53722 131172 53728
rect 131132 52601 131160 53722
rect 131212 53712 131264 53718
rect 131316 53689 131344 55082
rect 131212 53654 131264 53660
rect 131302 53680 131358 53689
rect 131224 53145 131252 53654
rect 131302 53615 131358 53624
rect 131210 53136 131266 53145
rect 131210 53071 131266 53080
rect 131118 52592 131174 52601
rect 131118 52527 131174 52536
rect 131212 52420 131264 52426
rect 131212 52362 131264 52368
rect 131224 51377 131252 52362
rect 131210 51368 131266 51377
rect 131210 51303 131266 51312
rect 131120 51060 131172 51066
rect 131120 51002 131172 51008
rect 131132 50289 131160 51002
rect 131212 50992 131264 50998
rect 131212 50934 131264 50940
rect 131224 50833 131252 50934
rect 131304 50924 131356 50930
rect 131304 50866 131356 50872
rect 131210 50824 131266 50833
rect 131210 50759 131266 50768
rect 131118 50280 131174 50289
rect 131118 50215 131174 50224
rect 131212 49700 131264 49706
rect 131212 49642 131264 49648
rect 131120 49632 131172 49638
rect 131120 49574 131172 49580
rect 131132 48521 131160 49574
rect 131224 49065 131252 49642
rect 131316 49609 131344 50866
rect 131302 49600 131358 49609
rect 131302 49535 131358 49544
rect 131210 49056 131266 49065
rect 131210 48991 131266 49000
rect 131118 48512 131174 48521
rect 131118 48447 131174 48456
rect 131212 48272 131264 48278
rect 131212 48214 131264 48220
rect 131224 47297 131252 48214
rect 131210 47288 131266 47297
rect 131210 47223 131266 47232
rect 131212 46912 131264 46918
rect 131212 46854 131264 46860
rect 131120 46844 131172 46850
rect 131120 46786 131172 46792
rect 131132 46209 131160 46786
rect 131224 46753 131252 46854
rect 131210 46744 131266 46753
rect 131210 46679 131266 46688
rect 131118 46200 131174 46209
rect 131118 46135 131174 46144
rect 131304 45552 131356 45558
rect 131304 45494 131356 45500
rect 131120 45484 131172 45490
rect 131120 45426 131172 45432
rect 131132 44985 131160 45426
rect 131212 45416 131264 45422
rect 131210 45384 131212 45393
rect 131264 45384 131266 45393
rect 131210 45319 131266 45328
rect 131118 44976 131174 44985
rect 131118 44911 131174 44920
rect 131316 44441 131344 45494
rect 131302 44432 131358 44441
rect 131302 44367 131358 44376
rect 131212 44124 131264 44130
rect 131212 44066 131264 44072
rect 131120 44056 131172 44062
rect 131120 43998 131172 44004
rect 131132 43217 131160 43998
rect 131224 43761 131252 44066
rect 131210 43752 131266 43761
rect 131210 43687 131266 43696
rect 131118 43208 131174 43217
rect 131118 43143 131174 43152
rect 131304 42832 131356 42838
rect 131304 42774 131356 42780
rect 131120 42764 131172 42770
rect 131120 42706 131172 42712
rect 131132 41993 131160 42706
rect 131212 42696 131264 42702
rect 131210 42664 131212 42673
rect 131264 42664 131266 42673
rect 131210 42599 131266 42608
rect 131118 41984 131174 41993
rect 131118 41919 131174 41928
rect 131120 41404 131172 41410
rect 131120 41346 131172 41352
rect 131132 40361 131160 41346
rect 131212 41336 131264 41342
rect 131212 41278 131264 41284
rect 131224 40905 131252 41278
rect 131210 40896 131266 40905
rect 131210 40831 131266 40840
rect 131118 40352 131174 40361
rect 131118 40287 131174 40296
rect 131212 38616 131264 38622
rect 131210 38584 131212 38593
rect 131264 38584 131266 38593
rect 131120 38548 131172 38554
rect 131210 38519 131266 38528
rect 131120 38490 131172 38496
rect 131132 37913 131160 38490
rect 131118 37904 131174 37913
rect 131118 37839 131174 37848
rect 131212 37256 131264 37262
rect 131212 37198 131264 37204
rect 131224 36145 131252 37198
rect 131316 36825 131344 42774
rect 131488 39364 131540 39370
rect 131488 39306 131540 39312
rect 131500 37369 131528 39306
rect 131486 37360 131542 37369
rect 131486 37295 131542 37304
rect 131302 36816 131358 36825
rect 131302 36751 131358 36760
rect 131210 36136 131266 36145
rect 131210 36071 131266 36080
rect 131212 35896 131264 35902
rect 131212 35838 131264 35844
rect 131120 35828 131172 35834
rect 131120 35770 131172 35776
rect 131132 35057 131160 35770
rect 131224 35601 131252 35838
rect 131210 35592 131266 35601
rect 131210 35527 131266 35536
rect 131118 35048 131174 35057
rect 131118 34983 131174 34992
rect 131120 33176 131172 33182
rect 131120 33118 131172 33124
rect 131132 32065 131160 33118
rect 131212 33108 131264 33114
rect 131212 33050 131264 33056
rect 131224 32745 131252 33050
rect 131210 32736 131266 32745
rect 131210 32671 131266 32680
rect 131118 32056 131174 32065
rect 131118 31991 131174 32000
rect 131212 31884 131264 31890
rect 131212 31826 131264 31832
rect 131224 31521 131252 31826
rect 131304 31816 131356 31822
rect 131304 31758 131356 31764
rect 131210 31512 131266 31521
rect 131210 31447 131266 31456
rect 131120 31068 131172 31074
rect 131120 31010 131172 31016
rect 131132 30433 131160 31010
rect 131316 30977 131344 31758
rect 131302 30968 131358 30977
rect 131302 30903 131358 30912
rect 131118 30424 131174 30433
rect 131118 30359 131174 30368
rect 131776 29306 131804 297298
rect 190472 267734 190500 304982
rect 190472 267706 190776 267734
rect 148324 260364 148376 260370
rect 148324 260306 148376 260312
rect 148336 252074 148364 260306
rect 153200 260296 153252 260302
rect 153200 260238 153252 260244
rect 148324 252068 148376 252074
rect 148324 252010 148376 252016
rect 153212 252006 153240 260238
rect 153200 252000 153252 252006
rect 153200 251942 153252 251948
rect 190748 249914 190776 267706
rect 193232 249914 193260 306342
rect 194600 282328 194652 282334
rect 194600 282270 194652 282276
rect 194612 267734 194640 282270
rect 197360 282260 197412 282266
rect 197360 282202 197412 282208
rect 197372 267734 197400 282202
rect 204272 267734 204300 325654
rect 207018 307184 207074 307193
rect 207018 307119 207074 307128
rect 207032 306406 207060 307119
rect 207020 306400 207072 306406
rect 207020 306342 207072 306348
rect 207018 305552 207074 305561
rect 207018 305487 207074 305496
rect 207032 305046 207060 305487
rect 207020 305040 207072 305046
rect 207020 304982 207072 304988
rect 208136 282402 208164 327383
rect 208124 282396 208176 282402
rect 208124 282338 208176 282344
rect 194612 267706 195376 267734
rect 197372 267706 197584 267734
rect 204272 267706 204576 267734
rect 195348 249914 195376 267706
rect 197556 249914 197584 267706
rect 202144 260296 202196 260302
rect 202144 260238 202196 260244
rect 201408 256148 201460 256154
rect 201408 256090 201460 256096
rect 201420 252550 201448 256090
rect 200396 252544 200448 252550
rect 200396 252486 200448 252492
rect 201408 252544 201460 252550
rect 201408 252486 201460 252492
rect 200408 249914 200436 252486
rect 190748 249886 191130 249914
rect 193232 249886 193430 249914
rect 195348 249886 195730 249914
rect 197556 249886 198030 249914
rect 200330 249886 200436 249914
rect 202156 249914 202184 260238
rect 204548 249914 204576 267706
rect 208228 253434 208256 331055
rect 208216 253428 208268 253434
rect 208216 253370 208268 253376
rect 207664 253292 207716 253298
rect 207664 253234 207716 253240
rect 207676 249914 207704 253234
rect 208320 253230 208348 332823
rect 209594 330032 209650 330041
rect 209594 329967 209650 329976
rect 209502 328536 209558 328545
rect 209502 328471 209558 328480
rect 209516 279682 209544 328471
rect 209608 280838 209636 329967
rect 209596 280832 209648 280838
rect 209596 280774 209648 280780
rect 209504 279676 209556 279682
rect 209504 279618 209556 279624
rect 209504 256216 209556 256222
rect 209504 256158 209556 256164
rect 208308 253224 208360 253230
rect 208308 253166 208360 253172
rect 202156 249886 202630 249914
rect 204548 249886 205022 249914
rect 207322 249886 207704 249914
rect 209516 249914 209544 256158
rect 209700 254794 209728 334047
rect 238574 299840 238630 299849
rect 238574 299775 238630 299784
rect 229098 298344 229154 298353
rect 227720 298308 227772 298314
rect 229098 298279 229154 298288
rect 227720 298250 227772 298256
rect 215852 298172 215904 298178
rect 215852 298114 215904 298120
rect 215864 298081 215892 298114
rect 227732 298081 227760 298250
rect 229112 298246 229140 298279
rect 229100 298240 229152 298246
rect 229100 298182 229152 298188
rect 215850 298072 215906 298081
rect 215850 298007 215906 298016
rect 224958 298072 225014 298081
rect 224958 298007 225014 298016
rect 226338 298072 226394 298081
rect 226338 298007 226394 298016
rect 227718 298072 227774 298081
rect 227718 298007 227774 298016
rect 213920 282396 213972 282402
rect 213920 282338 213972 282344
rect 211528 261724 211580 261730
rect 211528 261666 211580 261672
rect 209688 254788 209740 254794
rect 209688 254730 209740 254736
rect 211540 249914 211568 261666
rect 213932 249914 213960 282338
rect 224972 282334 225000 298007
rect 224960 282328 225012 282334
rect 224960 282270 225012 282276
rect 218060 280900 218112 280906
rect 218060 280842 218112 280848
rect 218072 267734 218100 280842
rect 222200 279676 222252 279682
rect 222200 279618 222252 279624
rect 222212 267734 222240 279618
rect 218072 267706 218560 267734
rect 222212 267706 223160 267734
rect 216128 260364 216180 260370
rect 216128 260306 216180 260312
rect 216140 249914 216168 260306
rect 218532 249914 218560 267706
rect 221464 256284 221516 256290
rect 221464 256226 221516 256232
rect 221476 249914 221504 256226
rect 209516 249886 209622 249914
rect 211540 249886 211922 249914
rect 213932 249886 214222 249914
rect 216140 249886 216522 249914
rect 218532 249886 218914 249914
rect 221214 249886 221504 249914
rect 223132 249914 223160 267706
rect 225328 260432 225380 260438
rect 225328 260374 225380 260380
rect 225340 249914 225368 260374
rect 226352 256154 226380 298007
rect 227732 256222 227760 298007
rect 229112 280906 229140 298182
rect 230478 298072 230534 298081
rect 230478 298007 230534 298016
rect 231950 298072 232006 298081
rect 231950 298007 232006 298016
rect 233238 298072 233294 298081
rect 233238 298007 233294 298016
rect 234710 298072 234766 298081
rect 234710 298007 234766 298016
rect 237194 298072 237250 298081
rect 237194 298007 237250 298016
rect 229282 297800 229338 297809
rect 229282 297735 229338 297744
rect 229296 297294 229324 297735
rect 229284 297288 229336 297294
rect 229284 297230 229336 297236
rect 229296 296714 229324 297230
rect 229204 296686 229324 296714
rect 229100 280900 229152 280906
rect 229100 280842 229152 280848
rect 229100 268184 229152 268190
rect 229100 268126 229152 268132
rect 227720 256216 227772 256222
rect 227720 256158 227772 256164
rect 226340 256148 226392 256154
rect 226340 256090 226392 256096
rect 228456 253904 228508 253910
rect 228456 253846 228508 253852
rect 228468 249914 228496 253846
rect 229112 250050 229140 268126
rect 229204 253910 229232 296686
rect 230492 260302 230520 298007
rect 231860 280832 231912 280838
rect 231860 280774 231912 280780
rect 230480 260296 230532 260302
rect 230480 260238 230532 260244
rect 231872 258074 231900 280774
rect 231964 261730 231992 298007
rect 231952 261724 232004 261730
rect 231952 261666 232004 261672
rect 231872 258046 232360 258074
rect 229192 253904 229244 253910
rect 229192 253846 229244 253852
rect 229112 250022 229968 250050
rect 223132 249886 223514 249914
rect 225340 249886 225814 249914
rect 228114 249886 228496 249914
rect 229940 249914 229968 250022
rect 232332 249914 232360 258046
rect 233252 256290 233280 298007
rect 234620 295996 234672 296002
rect 234620 295938 234672 295944
rect 234632 267734 234660 295938
rect 234724 268190 234752 298007
rect 234712 268184 234764 268190
rect 234712 268126 234764 268132
rect 234632 267706 234752 267734
rect 233240 256284 233292 256290
rect 233240 256226 233292 256232
rect 234724 249914 234752 267706
rect 237208 260302 237236 298007
rect 237378 297936 237434 297945
rect 237378 297871 237434 297880
rect 237286 297800 237342 297809
rect 237286 297735 237342 297744
rect 237196 260296 237248 260302
rect 237196 260238 237248 260244
rect 237300 252498 237328 297735
rect 237392 282266 237420 297871
rect 238588 297129 238616 299775
rect 243082 299704 243138 299713
rect 243082 299639 243138 299648
rect 238666 298072 238722 298081
rect 238666 298007 238722 298016
rect 240138 298072 240194 298081
rect 240138 298007 240194 298016
rect 241426 298072 241482 298081
rect 241426 298007 241482 298016
rect 242898 298072 242954 298081
rect 242898 298007 242954 298016
rect 238574 297120 238630 297129
rect 238574 297055 238630 297064
rect 237380 282260 237432 282266
rect 237380 282202 237432 282208
rect 237300 252470 237512 252498
rect 237484 249914 237512 252470
rect 238680 252210 238708 298007
rect 238758 297936 238814 297945
rect 238758 297871 238814 297880
rect 238772 253298 238800 297871
rect 240046 297120 240102 297129
rect 240046 297055 240102 297064
rect 239404 253428 239456 253434
rect 239404 253370 239456 253376
rect 238760 253292 238812 253298
rect 238760 253234 238812 253240
rect 238668 252204 238720 252210
rect 238668 252146 238720 252152
rect 229940 249886 230414 249914
rect 232332 249886 232806 249914
rect 234724 249886 235106 249914
rect 237406 249886 237512 249914
rect 239416 249914 239444 253370
rect 240060 253298 240088 297055
rect 240152 260370 240180 298007
rect 240140 260364 240192 260370
rect 240140 260306 240192 260312
rect 240048 253292 240100 253298
rect 240048 253234 240100 253240
rect 241440 252142 241468 298007
rect 241518 297936 241574 297945
rect 241518 297871 241574 297880
rect 241532 260438 241560 297871
rect 242806 297800 242862 297809
rect 242806 297735 242862 297744
rect 242820 268394 242848 297735
rect 242912 296002 242940 298007
rect 243096 297945 243124 299639
rect 244094 298072 244150 298081
rect 244094 298007 244150 298016
rect 244278 298072 244334 298081
rect 244278 298007 244334 298016
rect 245566 298072 245622 298081
rect 245566 298007 245622 298016
rect 246854 298072 246910 298081
rect 246854 298007 246910 298016
rect 248234 298072 248290 298081
rect 248234 298007 248290 298016
rect 249706 298072 249762 298081
rect 249706 298007 249762 298016
rect 250994 298072 251050 298081
rect 250994 298007 251050 298016
rect 252374 298072 252430 298081
rect 252374 298007 252430 298016
rect 253754 298072 253810 298081
rect 253754 298007 253810 298016
rect 255134 298072 255190 298081
rect 255134 298007 255190 298016
rect 256514 298072 256570 298081
rect 256514 298007 256570 298016
rect 257894 298072 257950 298081
rect 257894 298007 257950 298016
rect 259182 298072 259238 298081
rect 259182 298007 259238 298016
rect 260654 298072 260710 298081
rect 260654 298007 260710 298016
rect 262034 298072 262090 298081
rect 262034 298007 262090 298016
rect 263506 298072 263562 298081
rect 263506 298007 263562 298016
rect 266174 298072 266230 298081
rect 266174 298007 266230 298016
rect 273074 298072 273130 298081
rect 273074 298007 273130 298016
rect 274546 298072 274602 298081
rect 274546 298007 274602 298016
rect 275926 298072 275982 298081
rect 275926 298007 275982 298016
rect 277306 298072 277362 298081
rect 277306 298007 277362 298016
rect 243082 297936 243138 297945
rect 243082 297871 243138 297880
rect 242900 295996 242952 296002
rect 242900 295938 242952 295944
rect 242808 268388 242860 268394
rect 242808 268330 242860 268336
rect 241520 260432 241572 260438
rect 241520 260374 241572 260380
rect 241612 260092 241664 260098
rect 241612 260034 241664 260040
rect 241428 252136 241480 252142
rect 241428 252078 241480 252084
rect 241624 249914 241652 260034
rect 244108 259010 244136 298007
rect 244186 297936 244242 297945
rect 244186 297871 244242 297880
rect 244096 259004 244148 259010
rect 244096 258946 244148 258952
rect 244200 257582 244228 297871
rect 244292 260098 244320 298007
rect 245580 273970 245608 298007
rect 246762 297936 246818 297945
rect 246762 297871 246818 297880
rect 245568 273964 245620 273970
rect 245568 273906 245620 273912
rect 246776 271862 246804 297871
rect 246764 271856 246816 271862
rect 246764 271798 246816 271804
rect 246868 261730 246896 298007
rect 246946 297800 247002 297809
rect 246946 297735 247002 297744
rect 246856 261724 246908 261730
rect 246856 261666 246908 261672
rect 244372 260296 244424 260302
rect 244372 260238 244424 260244
rect 244280 260092 244332 260098
rect 244280 260034 244332 260040
rect 244188 257576 244240 257582
rect 244188 257518 244240 257524
rect 244384 249914 244412 260238
rect 246960 257718 246988 297735
rect 248248 280838 248276 298007
rect 248326 297936 248382 297945
rect 248326 297871 248382 297880
rect 249614 297936 249670 297945
rect 249614 297871 249670 297880
rect 248236 280832 248288 280838
rect 248236 280774 248288 280780
rect 248340 263158 248368 297871
rect 248420 271856 248472 271862
rect 248420 271798 248472 271804
rect 248432 267734 248460 271798
rect 248432 267706 248552 267734
rect 248328 263152 248380 263158
rect 248328 263094 248380 263100
rect 246948 257712 247000 257718
rect 246948 257654 247000 257660
rect 246396 253224 246448 253230
rect 246396 253166 246448 253172
rect 239416 249886 239706 249914
rect 241624 249886 242006 249914
rect 244306 249886 244412 249914
rect 246408 249914 246436 253166
rect 248524 249914 248552 267706
rect 249628 258942 249656 297871
rect 249616 258936 249668 258942
rect 249616 258878 249668 258884
rect 249720 253230 249748 298007
rect 251008 260302 251036 298007
rect 251086 297936 251142 297945
rect 251086 297871 251142 297880
rect 252282 297936 252338 297945
rect 252282 297871 252338 297880
rect 250996 260296 251048 260302
rect 250996 260238 251048 260244
rect 251100 258874 251128 297871
rect 252296 263090 252324 297871
rect 252284 263084 252336 263090
rect 252284 263026 252336 263032
rect 252388 263022 252416 298007
rect 252466 297800 252522 297809
rect 252466 297735 252522 297744
rect 252376 263016 252428 263022
rect 252376 262958 252428 262964
rect 252480 260506 252508 297735
rect 253768 264450 253796 298007
rect 253846 297936 253902 297945
rect 253846 297871 253902 297880
rect 253756 264444 253808 264450
rect 253756 264386 253808 264392
rect 252468 260500 252520 260506
rect 252468 260442 252520 260448
rect 253860 260438 253888 297871
rect 255148 264382 255176 298007
rect 255226 297936 255282 297945
rect 255226 297871 255282 297880
rect 255136 264376 255188 264382
rect 255136 264318 255188 264324
rect 255240 261866 255268 297871
rect 256528 264314 256556 298007
rect 256606 297936 256662 297945
rect 256606 297871 256662 297880
rect 257802 297936 257858 297945
rect 257802 297871 257858 297880
rect 256516 264308 256568 264314
rect 256516 264250 256568 264256
rect 255228 261860 255280 261866
rect 255228 261802 255280 261808
rect 256620 261798 256648 297871
rect 257816 265810 257844 297871
rect 257804 265804 257856 265810
rect 257804 265746 257856 265752
rect 256608 261792 256660 261798
rect 256608 261734 256660 261740
rect 255504 261724 255556 261730
rect 255504 261666 255556 261672
rect 253848 260432 253900 260438
rect 253848 260374 253900 260380
rect 251088 258868 251140 258874
rect 251088 258810 251140 258816
rect 253204 254788 253256 254794
rect 253204 254730 253256 254736
rect 249708 253224 249760 253230
rect 249708 253166 249760 253172
rect 251180 252204 251232 252210
rect 251180 252146 251232 252152
rect 251192 249914 251220 252146
rect 253216 249914 253244 254730
rect 255516 249914 255544 261666
rect 257908 256290 257936 298007
rect 257986 297800 258042 297809
rect 257986 297735 258042 297744
rect 257896 256284 257948 256290
rect 257896 256226 257948 256232
rect 258000 254794 258028 297735
rect 259196 265674 259224 298007
rect 259366 297936 259422 297945
rect 259366 297871 259422 297880
rect 259274 297800 259330 297809
rect 259274 297735 259330 297744
rect 259288 265742 259316 297735
rect 259276 265736 259328 265742
rect 259276 265678 259328 265684
rect 259184 265668 259236 265674
rect 259184 265610 259236 265616
rect 259380 261730 259408 297871
rect 259460 280832 259512 280838
rect 259460 280774 259512 280780
rect 259472 267734 259500 280774
rect 259472 267706 260144 267734
rect 259368 261724 259420 261730
rect 259368 261666 259420 261672
rect 257988 254788 258040 254794
rect 257988 254730 258040 254736
rect 258080 253292 258132 253298
rect 258080 253234 258132 253240
rect 258092 249914 258120 253234
rect 260116 249914 260144 267706
rect 260668 267170 260696 298007
rect 260746 297936 260802 297945
rect 260746 297871 260802 297880
rect 260656 267164 260708 267170
rect 260656 267106 260708 267112
rect 260760 257650 260788 297871
rect 262048 267102 262076 298007
rect 262126 297936 262182 297945
rect 262126 297871 262182 297880
rect 263414 297936 263470 297945
rect 263414 297871 263470 297880
rect 262036 267096 262088 267102
rect 262036 267038 262088 267044
rect 260748 257644 260800 257650
rect 260748 257586 260800 257592
rect 262140 256222 262168 297871
rect 263428 267034 263456 297871
rect 263416 267028 263468 267034
rect 263416 266970 263468 266976
rect 262128 256216 262180 256222
rect 262128 256158 262180 256164
rect 263520 256154 263548 298007
rect 264794 296984 264850 296993
rect 264794 296919 264850 296928
rect 264808 268462 264836 296919
rect 264886 296848 264942 296857
rect 264886 296783 264942 296792
rect 264796 268456 264848 268462
rect 264796 268398 264848 268404
rect 263508 256148 263560 256154
rect 263508 256090 263560 256096
rect 264900 253706 264928 296783
rect 266188 282334 266216 298007
rect 267646 297120 267702 297129
rect 267646 297055 267702 297064
rect 267462 296984 267518 296993
rect 267462 296919 267518 296928
rect 266266 296848 266322 296857
rect 266266 296783 266322 296792
rect 266176 282328 266228 282334
rect 266176 282270 266228 282276
rect 264888 253700 264940 253706
rect 264888 253642 264940 253648
rect 266280 253638 266308 296783
rect 267476 282266 267504 296919
rect 267554 296848 267610 296857
rect 267554 296783 267610 296792
rect 267464 282260 267516 282266
rect 267464 282202 267516 282208
rect 267568 268394 267596 296783
rect 266360 268388 266412 268394
rect 266360 268330 266412 268336
rect 267556 268388 267608 268394
rect 267556 268330 267608 268336
rect 266372 267734 266400 268330
rect 266372 267706 267136 267734
rect 266268 253632 266320 253638
rect 266268 253574 266320 253580
rect 264980 253224 265032 253230
rect 264980 253166 265032 253172
rect 262588 252136 262640 252142
rect 262588 252078 262640 252084
rect 262600 249914 262628 252078
rect 264992 249914 265020 253166
rect 267108 249914 267136 267706
rect 267660 253570 267688 297055
rect 269026 296848 269082 296857
rect 269026 296783 269082 296792
rect 270406 296848 270462 296857
rect 270406 296783 270462 296792
rect 271786 296848 271842 296857
rect 271786 296783 271842 296792
rect 267648 253564 267700 253570
rect 267648 253506 267700 253512
rect 269040 253502 269068 296783
rect 269304 260296 269356 260302
rect 269304 260238 269356 260244
rect 269028 253496 269080 253502
rect 269028 253438 269080 253444
rect 269316 249914 269344 260238
rect 270420 253434 270448 296783
rect 270408 253428 270460 253434
rect 270408 253370 270460 253376
rect 271800 253366 271828 296783
rect 273088 260370 273116 298007
rect 273166 296848 273222 296857
rect 273166 296783 273222 296792
rect 273076 260364 273128 260370
rect 273076 260306 273128 260312
rect 273180 260302 273208 296783
rect 274088 260500 274140 260506
rect 274088 260442 274140 260448
rect 273168 260296 273220 260302
rect 273168 260238 273220 260244
rect 271880 257576 271932 257582
rect 271880 257518 271932 257524
rect 271788 253360 271840 253366
rect 271788 253302 271840 253308
rect 271892 249914 271920 257518
rect 274100 249914 274128 260442
rect 274560 253298 274588 298007
rect 274548 253292 274600 253298
rect 274548 253234 274600 253240
rect 275940 253230 275968 298007
rect 276296 259004 276348 259010
rect 276296 258946 276348 258952
rect 275928 253224 275980 253230
rect 275928 253166 275980 253172
rect 276308 249914 276336 258946
rect 277320 257582 277348 298007
rect 341524 297220 341576 297226
rect 341524 297162 341576 297168
rect 280160 273964 280212 273970
rect 280160 273906 280212 273912
rect 280172 267734 280200 273906
rect 280172 267706 280936 267734
rect 278780 260432 278832 260438
rect 278780 260374 278832 260380
rect 277308 257576 277360 257582
rect 277308 257518 277360 257524
rect 278792 249914 278820 260374
rect 280908 249914 280936 267706
rect 341064 267164 341116 267170
rect 341064 267106 341116 267112
rect 327264 265804 327316 265810
rect 327264 265746 327316 265752
rect 313280 264444 313332 264450
rect 313280 264386 313332 264392
rect 290280 263152 290332 263158
rect 290280 263094 290332 263100
rect 283288 261860 283340 261866
rect 283288 261802 283340 261808
rect 283300 249914 283328 261802
rect 287888 261792 287940 261798
rect 287888 261734 287940 261740
rect 285680 257712 285732 257718
rect 285680 257654 285732 257660
rect 285692 249914 285720 257654
rect 287900 249914 287928 261734
rect 290292 249914 290320 263094
rect 304080 263084 304132 263090
rect 304080 263026 304132 263032
rect 302332 261724 302384 261730
rect 302332 261666 302384 261672
rect 294880 258936 294932 258942
rect 294880 258878 294932 258884
rect 292580 254788 292632 254794
rect 292580 254730 292632 254736
rect 292592 249914 292620 254730
rect 294892 249914 294920 258878
rect 299480 258868 299532 258874
rect 299480 258810 299532 258816
rect 297180 256284 297232 256290
rect 297180 256226 297232 256232
rect 297192 249914 297220 256226
rect 299492 249914 299520 258810
rect 302344 249914 302372 261666
rect 246408 249886 246698 249914
rect 248524 249886 248998 249914
rect 251192 249886 251298 249914
rect 253216 249886 253598 249914
rect 255516 249886 255898 249914
rect 258092 249886 258198 249914
rect 260116 249886 260590 249914
rect 262600 249886 262890 249914
rect 264992 249886 265190 249914
rect 267108 249886 267490 249914
rect 269316 249886 269790 249914
rect 271892 249886 272090 249914
rect 274100 249886 274482 249914
rect 276308 249886 276782 249914
rect 278792 249886 279082 249914
rect 280908 249886 281382 249914
rect 283300 249886 283682 249914
rect 285692 249886 285982 249914
rect 287900 249886 288374 249914
rect 290292 249886 290674 249914
rect 292592 249886 292974 249914
rect 294892 249886 295274 249914
rect 297192 249886 297574 249914
rect 299492 249886 299874 249914
rect 302266 249886 302372 249914
rect 304092 249914 304120 263026
rect 309232 263016 309284 263022
rect 309232 262958 309284 262964
rect 306564 257644 306616 257650
rect 306564 257586 306616 257592
rect 306576 249914 306604 257586
rect 309244 249914 309272 262958
rect 311164 256216 311216 256222
rect 311164 256158 311216 256164
rect 304092 249886 304566 249914
rect 306576 249886 306866 249914
rect 309166 249886 309272 249914
rect 311176 249914 311204 256158
rect 313292 249914 313320 264386
rect 318064 264376 318116 264382
rect 318064 264318 318116 264324
rect 316040 256148 316092 256154
rect 316040 256090 316092 256096
rect 316052 249914 316080 256090
rect 318076 249914 318104 264318
rect 322940 264308 322992 264314
rect 322940 264250 322992 264256
rect 320364 253700 320416 253706
rect 320364 253642 320416 253648
rect 320376 249914 320404 253642
rect 322952 249914 322980 264250
rect 324964 253632 325016 253638
rect 324964 253574 325016 253580
rect 324976 249914 325004 253574
rect 327276 249914 327304 265746
rect 331864 265736 331916 265742
rect 331864 265678 331916 265684
rect 329840 253564 329892 253570
rect 329840 253506 329892 253512
rect 329852 249914 329880 253506
rect 331876 249914 331904 265678
rect 336740 265668 336792 265674
rect 336740 265610 336792 265616
rect 334348 253496 334400 253502
rect 334348 253438 334400 253444
rect 334360 249914 334388 253438
rect 336752 249914 336780 265610
rect 338948 253428 339000 253434
rect 338948 253370 339000 253376
rect 338960 249914 338988 253370
rect 341076 249914 341104 267106
rect 341536 252142 341564 297162
rect 345664 297152 345716 297158
rect 345664 297094 345716 297100
rect 345572 267096 345624 267102
rect 345572 267038 345624 267044
rect 343640 253360 343692 253366
rect 343640 253302 343692 253308
rect 341524 252136 341576 252142
rect 341524 252078 341576 252084
rect 343652 249914 343680 253302
rect 345584 250050 345612 267038
rect 345676 252210 345704 297094
rect 409052 297084 409104 297090
rect 409052 297026 409104 297032
rect 408868 297016 408920 297022
rect 408868 296958 408920 296964
rect 371240 291848 371292 291854
rect 371240 291790 371292 291796
rect 358820 282328 358872 282334
rect 358820 282270 358872 282276
rect 354680 268456 354732 268462
rect 354680 268398 354732 268404
rect 354692 267734 354720 268398
rect 358832 267734 358860 282270
rect 364340 282260 364392 282266
rect 364340 282202 364392 282208
rect 354692 267706 355088 267734
rect 358832 267706 359688 267734
rect 350540 267028 350592 267034
rect 350540 266970 350592 266976
rect 348056 260364 348108 260370
rect 348056 260306 348108 260312
rect 345664 252204 345716 252210
rect 345664 252146 345716 252152
rect 345584 250022 345888 250050
rect 345860 249914 345888 250022
rect 348068 249914 348096 260306
rect 350552 249914 350580 266970
rect 352656 260296 352708 260302
rect 352656 260238 352708 260244
rect 352668 249914 352696 260238
rect 355060 249914 355088 267706
rect 357532 253292 357584 253298
rect 357532 253234 357584 253240
rect 357544 249914 357572 253234
rect 359660 249914 359688 267706
rect 362132 253224 362184 253230
rect 362132 253166 362184 253172
rect 362144 249914 362172 253166
rect 364352 249914 364380 282202
rect 368480 268388 368532 268394
rect 368480 268330 368532 268336
rect 368492 267734 368520 268330
rect 368492 267706 368888 267734
rect 366732 257576 366784 257582
rect 366732 257518 366784 257524
rect 366744 249914 366772 257518
rect 368860 249914 368888 267706
rect 371252 249914 371280 291790
rect 389180 279608 389232 279614
rect 389180 279550 389232 279556
rect 374000 279540 374052 279546
rect 374000 279482 374052 279488
rect 374012 267734 374040 279482
rect 389192 267734 389220 279550
rect 374012 267706 374132 267734
rect 389192 267706 389864 267734
rect 374104 249914 374132 267706
rect 387800 261656 387852 261662
rect 387800 261598 387852 261604
rect 375932 257372 375984 257378
rect 375932 257314 375984 257320
rect 311176 249886 311466 249914
rect 313292 249886 313766 249914
rect 316052 249886 316158 249914
rect 318076 249886 318458 249914
rect 320376 249886 320758 249914
rect 322952 249886 323058 249914
rect 324976 249886 325358 249914
rect 327276 249886 327658 249914
rect 329852 249886 330050 249914
rect 331876 249886 332350 249914
rect 334360 249886 334650 249914
rect 336752 249886 336950 249914
rect 338960 249886 339250 249914
rect 341076 249886 341550 249914
rect 343652 249886 343942 249914
rect 345860 249886 346242 249914
rect 348068 249886 348542 249914
rect 350552 249886 350842 249914
rect 352668 249886 353142 249914
rect 355060 249886 355442 249914
rect 357544 249886 357834 249914
rect 359660 249886 360134 249914
rect 362144 249886 362434 249914
rect 364352 249886 364734 249914
rect 366744 249886 367034 249914
rect 368860 249886 369334 249914
rect 371252 249886 371726 249914
rect 374026 249886 374132 249914
rect 375944 249914 375972 257314
rect 378324 252068 378376 252074
rect 378324 252010 378376 252016
rect 378336 249914 378364 252010
rect 385316 252000 385368 252006
rect 385316 251942 385368 251948
rect 380992 251932 381044 251938
rect 380992 251874 381044 251880
rect 381004 249914 381032 251874
rect 382924 251864 382976 251870
rect 382924 251806 382976 251812
rect 375944 249886 376326 249914
rect 378336 249886 378626 249914
rect 380926 249886 381032 249914
rect 382936 249914 382964 251806
rect 385328 249914 385356 251942
rect 387812 249914 387840 261598
rect 389836 249914 389864 267706
rect 399024 264240 399076 264246
rect 399024 264182 399076 264188
rect 392032 261588 392084 261594
rect 392032 261530 392084 261536
rect 392044 249914 392072 261530
rect 396724 257508 396776 257514
rect 396724 257450 396776 257456
rect 394700 257440 394752 257446
rect 394700 257382 394752 257388
rect 394712 249914 394740 257382
rect 396736 249914 396764 257450
rect 399036 249914 399064 264182
rect 403624 260228 403676 260234
rect 403624 260170 403676 260176
rect 401600 260160 401652 260166
rect 401600 260102 401652 260108
rect 401612 249914 401640 260102
rect 403636 249914 403664 260170
rect 408500 252204 408552 252210
rect 408500 252146 408552 252152
rect 406108 252136 406160 252142
rect 406108 252078 406160 252084
rect 406120 249914 406148 252078
rect 408512 249914 408540 252146
rect 382936 249886 383226 249914
rect 385328 249886 385618 249914
rect 387812 249886 387918 249914
rect 389836 249886 390218 249914
rect 392044 249886 392518 249914
rect 394712 249886 394818 249914
rect 396736 249886 397118 249914
rect 399036 249886 399510 249914
rect 401612 249886 401810 249914
rect 403636 249886 404110 249914
rect 406120 249886 406410 249914
rect 408512 249886 408710 249914
rect 186320 249756 186372 249762
rect 186320 249698 186372 249704
rect 186332 249529 186360 249698
rect 408880 249665 408908 296958
rect 408960 296744 409012 296750
rect 408960 296686 409012 296692
rect 408972 251841 409000 296686
rect 408958 251832 409014 251841
rect 408958 251767 409014 251776
rect 408866 249656 408922 249665
rect 408866 249591 408922 249600
rect 186318 249520 186374 249529
rect 186318 249455 186374 249464
rect 186412 248396 186464 248402
rect 186412 248338 186464 248344
rect 186320 248328 186372 248334
rect 186318 248296 186320 248305
rect 186372 248296 186374 248305
rect 186318 248231 186374 248240
rect 186424 247217 186452 248338
rect 186410 247208 186466 247217
rect 186410 247143 186466 247152
rect 186320 247036 186372 247042
rect 186320 246978 186372 246984
rect 186332 245993 186360 246978
rect 187148 246356 187200 246362
rect 187148 246298 187200 246304
rect 186318 245984 186374 245993
rect 186318 245919 186374 245928
rect 186320 245608 186372 245614
rect 186320 245550 186372 245556
rect 186332 244905 186360 245550
rect 186318 244896 186374 244905
rect 186318 244831 186374 244840
rect 186320 244248 186372 244254
rect 186320 244190 186372 244196
rect 186332 243681 186360 244190
rect 186318 243672 186374 243681
rect 186318 243607 186374 243616
rect 186320 242888 186372 242894
rect 186320 242830 186372 242836
rect 186332 242593 186360 242830
rect 186318 242584 186374 242593
rect 186318 242519 186374 242528
rect 186320 241460 186372 241466
rect 186320 241402 186372 241408
rect 186332 241369 186360 241402
rect 186318 241360 186374 241369
rect 186318 241295 186374 241304
rect 186318 240136 186374 240145
rect 186318 240071 186374 240080
rect 186412 240100 186464 240106
rect 186332 240038 186360 240071
rect 186412 240042 186464 240048
rect 186320 240032 186372 240038
rect 186320 239974 186372 239980
rect 186424 239057 186452 240042
rect 186410 239048 186466 239057
rect 186410 238983 186466 238992
rect 187160 237833 187188 246298
rect 409064 241618 409092 297026
rect 409328 296948 409380 296954
rect 409328 296890 409380 296896
rect 409236 296880 409288 296886
rect 409236 296822 409288 296828
rect 409144 296812 409196 296818
rect 409144 296754 409196 296760
rect 409156 243658 409184 296754
rect 409248 245562 409276 296822
rect 409340 247761 409368 296890
rect 409972 287700 410024 287706
rect 409972 287642 410024 287648
rect 409880 279472 409932 279478
rect 409880 279414 409932 279420
rect 409418 248296 409474 248305
rect 409418 248231 409474 248240
rect 409326 247752 409382 247761
rect 409326 247687 409382 247696
rect 409326 245576 409382 245585
rect 409248 245534 409326 245562
rect 409326 245511 409382 245520
rect 409326 243672 409382 243681
rect 409156 243630 409326 243658
rect 409326 243607 409382 243616
rect 409326 241632 409382 241641
rect 409064 241590 409326 241618
rect 409326 241567 409382 241576
rect 409432 238754 409460 248231
rect 408880 238726 409460 238754
rect 187146 237824 187202 237833
rect 187146 237759 187202 237768
rect 186320 237380 186372 237386
rect 186320 237322 186372 237328
rect 186332 236745 186360 237322
rect 186318 236736 186374 236745
rect 186318 236671 186374 236680
rect 186320 235952 186372 235958
rect 186320 235894 186372 235900
rect 186332 235521 186360 235894
rect 186318 235512 186374 235521
rect 186318 235447 186374 235456
rect 186320 234592 186372 234598
rect 186320 234534 186372 234540
rect 186332 234433 186360 234534
rect 186318 234424 186374 234433
rect 186318 234359 186374 234368
rect 186412 233232 186464 233238
rect 186318 233200 186374 233209
rect 186412 233174 186464 233180
rect 186318 233135 186320 233144
rect 186372 233135 186374 233144
rect 186320 233106 186372 233112
rect 186424 232121 186452 233174
rect 186410 232112 186466 232121
rect 186410 232047 186466 232056
rect 186320 231804 186372 231810
rect 186320 231746 186372 231752
rect 186332 230897 186360 231746
rect 186318 230888 186374 230897
rect 186318 230823 186374 230832
rect 186320 230444 186372 230450
rect 186320 230386 186372 230392
rect 186332 229673 186360 230386
rect 186318 229664 186374 229673
rect 186318 229599 186374 229608
rect 408880 229094 408908 238726
rect 408880 229066 409368 229094
rect 186318 228576 186374 228585
rect 186318 228511 186374 228520
rect 186332 227798 186360 228511
rect 169024 227792 169076 227798
rect 169024 227734 169076 227740
rect 186320 227792 186372 227798
rect 186320 227734 186372 227740
rect 148324 226364 148376 226370
rect 148324 226306 148376 226312
rect 133236 225004 133288 225010
rect 133236 224946 133288 224952
rect 131856 169788 131908 169794
rect 131856 169730 131908 169736
rect 131868 100473 131896 169730
rect 133144 130552 133196 130558
rect 133144 130494 133196 130500
rect 132040 128308 132092 128314
rect 132040 128250 132092 128256
rect 132052 127401 132080 128250
rect 132224 128240 132276 128246
rect 132224 128182 132276 128188
rect 132236 127945 132264 128182
rect 132222 127936 132278 127945
rect 132222 127871 132278 127880
rect 132038 127392 132094 127401
rect 132038 127327 132094 127336
rect 132040 126880 132092 126886
rect 132040 126822 132092 126828
rect 132052 125633 132080 126822
rect 132038 125624 132094 125633
rect 132038 125559 132094 125568
rect 132224 124160 132276 124166
rect 132224 124102 132276 124108
rect 132236 123865 132264 124102
rect 132222 123856 132278 123865
rect 132222 123791 132278 123800
rect 131948 121440 132000 121446
rect 131948 121382 132000 121388
rect 131960 120329 131988 121382
rect 131946 120320 132002 120329
rect 131946 120255 132002 120264
rect 132224 120080 132276 120086
rect 132224 120022 132276 120028
rect 132236 119785 132264 120022
rect 132222 119776 132278 119785
rect 132222 119711 132278 119720
rect 132132 111784 132184 111790
rect 132132 111726 132184 111732
rect 132144 111625 132172 111726
rect 132130 111616 132186 111625
rect 132130 111551 132186 111560
rect 131854 100464 131910 100473
rect 131854 100399 131910 100408
rect 131856 98048 131908 98054
rect 131856 97990 131908 97996
rect 131868 64297 131896 97990
rect 132224 96008 132276 96014
rect 132224 95950 132276 95956
rect 132236 95305 132264 95950
rect 132222 95296 132278 95305
rect 132222 95231 132278 95240
rect 131948 93900 132000 93906
rect 131948 93842 132000 93848
rect 131854 64288 131910 64297
rect 131854 64223 131910 64232
rect 131960 62529 131988 93842
rect 132224 89616 132276 89622
rect 132224 89558 132276 89564
rect 132236 89457 132264 89558
rect 132222 89448 132278 89457
rect 132222 89383 132278 89392
rect 132040 87032 132092 87038
rect 132040 86974 132092 86980
rect 131946 62520 132002 62529
rect 131946 62455 132002 62464
rect 132052 58993 132080 86974
rect 132224 85536 132276 85542
rect 132224 85478 132276 85484
rect 132236 85377 132264 85478
rect 132222 85368 132278 85377
rect 132222 85303 132278 85312
rect 132224 84856 132276 84862
rect 132224 84798 132276 84804
rect 132236 84153 132264 84798
rect 132222 84144 132278 84153
rect 132222 84079 132278 84088
rect 132224 81388 132276 81394
rect 132224 81330 132276 81336
rect 132236 81161 132264 81330
rect 132222 81152 132278 81161
rect 132222 81087 132278 81096
rect 132500 75200 132552 75206
rect 132500 75142 132552 75148
rect 132316 73228 132368 73234
rect 132316 73170 132368 73176
rect 132224 63504 132276 63510
rect 132224 63446 132276 63452
rect 132236 63073 132264 63446
rect 132222 63064 132278 63073
rect 132222 62999 132278 63008
rect 132132 62008 132184 62014
rect 132132 61950 132184 61956
rect 132144 61305 132172 61950
rect 132130 61296 132186 61305
rect 132130 61231 132186 61240
rect 132224 60648 132276 60654
rect 132224 60590 132276 60596
rect 132236 60217 132264 60590
rect 132222 60208 132278 60217
rect 132222 60143 132278 60152
rect 132038 58984 132094 58993
rect 132038 58919 132094 58928
rect 132224 56568 132276 56574
rect 132224 56510 132276 56516
rect 132236 56137 132264 56510
rect 132222 56128 132278 56137
rect 132222 56063 132278 56072
rect 131856 52488 131908 52494
rect 131856 52430 131908 52436
rect 131868 41449 131896 52430
rect 132328 52057 132356 73170
rect 132512 71913 132540 75142
rect 132498 71904 132554 71913
rect 132498 71839 132554 71848
rect 132500 55888 132552 55894
rect 132500 55830 132552 55836
rect 132512 54369 132540 55830
rect 132498 54360 132554 54369
rect 132498 54295 132554 54304
rect 132314 52048 132370 52057
rect 132314 51983 132370 51992
rect 132040 48340 132092 48346
rect 132040 48282 132092 48288
rect 131948 48068 132000 48074
rect 131948 48010 132000 48016
rect 131960 47841 131988 48010
rect 131946 47832 132002 47841
rect 131946 47767 132002 47776
rect 132052 45554 132080 48282
rect 132500 46980 132552 46986
rect 132500 46922 132552 46928
rect 131960 45526 132080 45554
rect 131854 41440 131910 41449
rect 131854 41375 131910 41384
rect 131960 39681 131988 45526
rect 131946 39672 132002 39681
rect 131946 39607 132002 39616
rect 132512 39137 132540 46922
rect 132498 39128 132554 39137
rect 132498 39063 132554 39072
rect 131856 38684 131908 38690
rect 131856 38626 131908 38632
rect 131868 34513 131896 38626
rect 132132 37324 132184 37330
rect 132132 37266 132184 37272
rect 131854 34504 131910 34513
rect 131854 34439 131910 34448
rect 132144 33833 132172 37266
rect 132224 35964 132276 35970
rect 132224 35906 132276 35912
rect 132130 33824 132186 33833
rect 132130 33759 132186 33768
rect 132236 33289 132264 35906
rect 132222 33280 132278 33289
rect 132222 33215 132278 33224
rect 131764 29300 131816 29306
rect 131764 29242 131816 29248
rect 130476 29096 130528 29102
rect 130476 29038 130528 29044
rect 79968 28960 80020 28966
rect 79968 28902 80020 28908
rect 133156 28354 133184 130494
rect 133248 128246 133276 224946
rect 145564 222216 145616 222222
rect 145564 222158 145616 222164
rect 135904 218068 135956 218074
rect 135904 218010 135956 218016
rect 134616 202904 134668 202910
rect 134616 202846 134668 202852
rect 134524 201544 134576 201550
rect 134524 201486 134576 201492
rect 133328 187740 133380 187746
rect 133328 187682 133380 187688
rect 133236 128240 133288 128246
rect 133236 128182 133288 128188
rect 133340 110430 133368 187682
rect 133512 158772 133564 158778
rect 133512 158714 133564 158720
rect 133420 157412 133472 157418
rect 133420 157354 133472 157360
rect 133328 110424 133380 110430
rect 133328 110366 133380 110372
rect 133432 95130 133460 157354
rect 133524 96014 133552 158714
rect 133604 154624 133656 154630
rect 133604 154566 133656 154572
rect 133512 96008 133564 96014
rect 133512 95950 133564 95956
rect 133420 95124 133472 95130
rect 133420 95066 133472 95072
rect 133616 93770 133644 154566
rect 134536 117230 134564 201486
rect 134628 118522 134656 202846
rect 134708 198756 134760 198762
rect 134708 198698 134760 198704
rect 134616 118516 134668 118522
rect 134616 118458 134668 118464
rect 134524 117224 134576 117230
rect 134524 117166 134576 117172
rect 134720 115530 134748 198698
rect 134800 161492 134852 161498
rect 134800 161434 134852 161440
rect 134708 115524 134760 115530
rect 134708 115466 134760 115472
rect 134524 110492 134576 110498
rect 134524 110434 134576 110440
rect 133696 101448 133748 101454
rect 133696 101390 133748 101396
rect 133604 93764 133656 93770
rect 133604 93706 133656 93712
rect 133236 92540 133288 92546
rect 133236 92482 133288 92488
rect 133248 62082 133276 92482
rect 133328 89752 133380 89758
rect 133328 89694 133380 89700
rect 133236 62076 133288 62082
rect 133236 62018 133288 62024
rect 133340 60654 133368 89694
rect 133420 85604 133472 85610
rect 133420 85546 133472 85552
rect 133328 60648 133380 60654
rect 133328 60590 133380 60596
rect 133432 59362 133460 85546
rect 133708 73166 133736 101390
rect 133696 73160 133748 73166
rect 133696 73102 133748 73108
rect 134536 71670 134564 110434
rect 134616 103556 134668 103562
rect 134616 103498 134668 103504
rect 134524 71664 134576 71670
rect 134524 71606 134576 71612
rect 133512 70440 133564 70446
rect 133512 70382 133564 70388
rect 133420 59356 133472 59362
rect 133420 59298 133472 59304
rect 133236 57996 133288 58002
rect 133236 57938 133288 57944
rect 133248 45558 133276 57938
rect 133328 53848 133380 53854
rect 133328 53790 133380 53796
rect 133236 45552 133288 45558
rect 133236 45494 133288 45500
rect 133340 42702 133368 53790
rect 133420 51128 133472 51134
rect 133420 51070 133472 51076
rect 133328 42696 133380 42702
rect 133328 42638 133380 42644
rect 133432 41342 133460 51070
rect 133524 50998 133552 70382
rect 134524 69080 134576 69086
rect 134524 69022 134576 69028
rect 133512 50992 133564 50998
rect 133512 50934 133564 50940
rect 134536 50930 134564 69022
rect 134628 67386 134656 103498
rect 134708 100768 134760 100774
rect 134708 100710 134760 100716
rect 134616 67380 134668 67386
rect 134616 67322 134668 67328
rect 134720 66162 134748 100710
rect 134812 96490 134840 161434
rect 135916 125526 135944 218010
rect 142804 215348 142856 215354
rect 142804 215290 142856 215296
rect 135996 212560 136048 212566
rect 135996 212502 136048 212508
rect 135904 125520 135956 125526
rect 135904 125462 135956 125468
rect 136008 122670 136036 212502
rect 140044 204332 140096 204338
rect 140044 204274 140096 204280
rect 137284 193248 137336 193254
rect 137284 193190 137336 193196
rect 136088 155984 136140 155990
rect 136088 155926 136140 155932
rect 135996 122664 136048 122670
rect 135996 122606 136048 122612
rect 135904 118720 135956 118726
rect 135904 118662 135956 118668
rect 134800 96484 134852 96490
rect 134800 96426 134852 96432
rect 134800 75948 134852 75954
rect 134800 75890 134852 75896
rect 134708 66156 134760 66162
rect 134708 66098 134760 66104
rect 134616 64932 134668 64938
rect 134616 64874 134668 64880
rect 134524 50924 134576 50930
rect 134524 50866 134576 50872
rect 134628 48074 134656 64874
rect 134708 60784 134760 60790
rect 134708 60726 134760 60732
rect 134616 48068 134668 48074
rect 134616 48010 134668 48016
rect 134720 46850 134748 60726
rect 134812 55146 134840 75890
rect 135916 75818 135944 118662
rect 136100 93838 136128 155926
rect 137296 113082 137324 193190
rect 137376 186380 137428 186386
rect 137376 186322 137428 186328
rect 137284 113076 137336 113082
rect 137284 113018 137336 113024
rect 137388 108934 137416 186322
rect 137468 179444 137520 179450
rect 137468 179386 137520 179392
rect 137376 108928 137428 108934
rect 137376 108870 137428 108876
rect 137480 106214 137508 179386
rect 138664 176724 138716 176730
rect 138664 176666 138716 176672
rect 137560 171148 137612 171154
rect 137560 171090 137612 171096
rect 137468 106208 137520 106214
rect 137468 106150 137520 106156
rect 137572 102066 137600 171090
rect 138676 104786 138704 176666
rect 138756 172576 138808 172582
rect 138756 172518 138808 172524
rect 138664 104780 138716 104786
rect 138664 104722 138716 104728
rect 138768 103358 138796 172518
rect 138848 153264 138900 153270
rect 138848 153206 138900 153212
rect 138756 103352 138808 103358
rect 138756 103294 138808 103300
rect 137560 102060 137612 102066
rect 137560 102002 137612 102008
rect 136088 93832 136140 93838
rect 136088 93774 136140 93780
rect 138860 92342 138888 153206
rect 140056 118590 140084 204274
rect 141424 194608 141476 194614
rect 141424 194550 141476 194556
rect 140136 190528 140188 190534
rect 140136 190470 140188 190476
rect 140044 118584 140096 118590
rect 140044 118526 140096 118532
rect 140148 111722 140176 190470
rect 140228 183592 140280 183598
rect 140228 183534 140280 183540
rect 140136 111716 140188 111722
rect 140136 111658 140188 111664
rect 140240 107506 140268 183534
rect 140320 180872 140372 180878
rect 140320 180814 140372 180820
rect 140332 107574 140360 180814
rect 141436 114374 141464 194550
rect 141516 184952 141568 184958
rect 141516 184894 141568 184900
rect 141424 114368 141476 114374
rect 141424 114310 141476 114316
rect 141424 109064 141476 109070
rect 141424 109006 141476 109012
rect 140320 107568 140372 107574
rect 140320 107510 140372 107516
rect 140228 107500 140280 107506
rect 140228 107442 140280 107448
rect 140044 106344 140096 106350
rect 140044 106286 140096 106292
rect 138848 92336 138900 92342
rect 138848 92278 138900 92284
rect 138664 88392 138716 88398
rect 138664 88334 138716 88340
rect 135996 82884 136048 82890
rect 135996 82826 136048 82832
rect 135904 75812 135956 75818
rect 135904 75754 135956 75760
rect 136008 57798 136036 82826
rect 136088 80096 136140 80102
rect 136088 80038 136140 80044
rect 135996 57792 136048 57798
rect 135996 57734 136048 57740
rect 136100 56506 136128 80038
rect 138676 60722 138704 88334
rect 138756 78736 138808 78742
rect 138756 78678 138808 78684
rect 138664 60716 138716 60722
rect 138664 60658 138716 60664
rect 136088 56500 136140 56506
rect 136088 56442 136140 56448
rect 138768 55214 138796 78678
rect 138848 76016 138900 76022
rect 138848 75958 138900 75964
rect 138756 55208 138808 55214
rect 138756 55150 138808 55156
rect 134800 55140 134852 55146
rect 134800 55082 134852 55088
rect 138860 53718 138888 75958
rect 140056 68882 140084 106286
rect 140136 102196 140188 102202
rect 140136 102138 140188 102144
rect 140044 68876 140096 68882
rect 140044 68818 140096 68824
rect 140148 67590 140176 102138
rect 140228 96688 140280 96694
rect 140228 96630 140280 96636
rect 140136 67584 140188 67590
rect 140136 67526 140188 67532
rect 140240 64802 140268 96630
rect 140320 95260 140372 95266
rect 140320 95202 140372 95208
rect 140228 64796 140280 64802
rect 140228 64738 140280 64744
rect 140332 63510 140360 95202
rect 141436 70310 141464 109006
rect 141528 109002 141556 184894
rect 141608 175296 141660 175302
rect 141608 175238 141660 175244
rect 141516 108996 141568 109002
rect 141516 108938 141568 108944
rect 141516 104916 141568 104922
rect 141516 104858 141568 104864
rect 141424 70304 141476 70310
rect 141424 70246 141476 70252
rect 141528 68950 141556 104858
rect 141620 103426 141648 175238
rect 141700 151836 141752 151842
rect 141700 151778 141752 151784
rect 141608 103420 141660 103426
rect 141608 103362 141660 103368
rect 141608 98116 141660 98122
rect 141608 98058 141660 98064
rect 141516 68944 141568 68950
rect 141516 68886 141568 68892
rect 141620 64870 141648 98058
rect 141712 92410 141740 151778
rect 142816 124098 142844 215290
rect 144184 200184 144236 200190
rect 144184 200126 144236 200132
rect 142896 136672 142948 136678
rect 142896 136614 142948 136620
rect 142804 124092 142856 124098
rect 142804 124034 142856 124040
rect 142804 120148 142856 120154
rect 142804 120090 142856 120096
rect 141792 116000 141844 116006
rect 141792 115942 141844 115948
rect 141700 92404 141752 92410
rect 141700 92346 141752 92352
rect 141804 74458 141832 115942
rect 142816 75886 142844 120090
rect 142908 84862 142936 136614
rect 142988 129804 143040 129810
rect 142988 129746 143040 129752
rect 142896 84856 142948 84862
rect 142896 84798 142948 84804
rect 142896 82952 142948 82958
rect 142896 82894 142948 82900
rect 142804 75880 142856 75886
rect 142804 75822 142856 75828
rect 141792 74452 141844 74458
rect 141792 74394 141844 74400
rect 141608 64864 141660 64870
rect 141608 64806 141660 64812
rect 140320 63504 140372 63510
rect 140320 63446 140372 63452
rect 142804 62144 142856 62150
rect 142804 62086 142856 62092
rect 141424 59424 141476 59430
rect 141424 59366 141476 59372
rect 140044 55276 140096 55282
rect 140044 55218 140096 55224
rect 138848 53712 138900 53718
rect 138848 53654 138900 53660
rect 134708 46844 134760 46850
rect 134708 46786 134760 46792
rect 140056 44062 140084 55218
rect 141436 45490 141464 59366
rect 142816 46918 142844 62086
rect 142908 57866 142936 82894
rect 143000 81326 143028 129746
rect 143080 127016 143132 127022
rect 143080 126958 143132 126964
rect 142988 81320 143040 81326
rect 142988 81262 143040 81268
rect 143092 79898 143120 126958
rect 144196 115938 144224 200126
rect 144276 178084 144328 178090
rect 144276 178026 144328 178032
rect 144184 115932 144236 115938
rect 144184 115874 144236 115880
rect 144288 104854 144316 178026
rect 144368 147688 144420 147694
rect 144368 147630 144420 147636
rect 144276 104848 144328 104854
rect 144276 104790 144328 104796
rect 144184 99408 144236 99414
rect 144184 99350 144236 99356
rect 143080 79892 143132 79898
rect 143080 79834 143132 79840
rect 144196 66230 144224 99350
rect 144380 89622 144408 147630
rect 144460 143608 144512 143614
rect 144460 143550 144512 143556
rect 144368 89616 144420 89622
rect 144368 89558 144420 89564
rect 144472 89010 144500 143550
rect 145576 126818 145604 222158
rect 145656 219496 145708 219502
rect 145656 219438 145708 219444
rect 145668 126886 145696 219438
rect 145748 211200 145800 211206
rect 145748 211142 145800 211148
rect 145656 126880 145708 126886
rect 145656 126822 145708 126828
rect 145564 126812 145616 126818
rect 145564 126754 145616 126760
rect 145564 124228 145616 124234
rect 145564 124170 145616 124176
rect 144460 89004 144512 89010
rect 144460 88946 144512 88952
rect 145576 78606 145604 124170
rect 145760 122738 145788 211142
rect 146944 202972 146996 202978
rect 146944 202914 146996 202920
rect 145748 122732 145800 122738
rect 145748 122674 145800 122680
rect 145748 120216 145800 120222
rect 145748 120158 145800 120164
rect 145656 117360 145708 117366
rect 145656 117302 145708 117308
rect 145564 78600 145616 78606
rect 145564 78542 145616 78548
rect 145668 74526 145696 117302
rect 145760 77178 145788 120158
rect 146956 117298 146984 202914
rect 147036 194676 147088 194682
rect 147036 194618 147088 194624
rect 146944 117292 146996 117298
rect 146944 117234 146996 117240
rect 147048 113150 147076 194618
rect 147128 191888 147180 191894
rect 147128 191830 147180 191836
rect 147036 113144 147088 113150
rect 147036 113086 147088 113092
rect 146944 111852 146996 111858
rect 146944 111794 146996 111800
rect 145748 77172 145800 77178
rect 145748 77114 145800 77120
rect 145656 74520 145708 74526
rect 145656 74462 145708 74468
rect 146956 71738 146984 111794
rect 147140 111790 147168 191830
rect 148336 129606 148364 226306
rect 157984 225072 158036 225078
rect 157984 225014 158036 225020
rect 151084 223644 151136 223650
rect 151084 223586 151136 223592
rect 149704 216708 149756 216714
rect 149704 216650 149756 216656
rect 148416 142180 148468 142186
rect 148416 142122 148468 142128
rect 148324 129600 148376 129606
rect 148324 129542 148376 129548
rect 147220 128376 147272 128382
rect 147220 128318 147272 128324
rect 147128 111784 147180 111790
rect 147128 111726 147180 111732
rect 147036 107704 147088 107710
rect 147036 107646 147088 107652
rect 146944 71732 146996 71738
rect 146944 71674 146996 71680
rect 147048 70378 147076 107646
rect 147128 106412 147180 106418
rect 147128 106354 147180 106360
rect 147036 70372 147088 70378
rect 147036 70314 147088 70320
rect 146944 69148 146996 69154
rect 146944 69090 146996 69096
rect 144276 66292 144328 66298
rect 144276 66234 144328 66240
rect 144184 66224 144236 66230
rect 144184 66166 144236 66172
rect 142896 57860 142948 57866
rect 142896 57802 142948 57808
rect 144288 49638 144316 66234
rect 146956 51066 146984 69090
rect 147140 69018 147168 106354
rect 147232 79966 147260 128318
rect 148428 86902 148456 142122
rect 148508 138032 148560 138038
rect 148508 137974 148560 137980
rect 148416 86896 148468 86902
rect 148416 86838 148468 86844
rect 148520 85474 148548 137974
rect 148600 135312 148652 135318
rect 148600 135254 148652 135260
rect 148508 85468 148560 85474
rect 148508 85410 148560 85416
rect 148612 84114 148640 135254
rect 148692 131164 148744 131170
rect 148692 131106 148744 131112
rect 148600 84108 148652 84114
rect 148600 84050 148652 84056
rect 148704 81394 148732 131106
rect 149716 124166 149744 216650
rect 149796 209840 149848 209846
rect 149796 209782 149848 209788
rect 149704 124160 149756 124166
rect 149704 124102 149756 124108
rect 149704 121508 149756 121514
rect 149704 121450 149756 121456
rect 148692 81388 148744 81394
rect 148692 81330 148744 81336
rect 147220 79960 147272 79966
rect 147220 79902 147272 79908
rect 149716 77246 149744 121450
rect 149808 121378 149836 209782
rect 151096 128314 151124 223586
rect 156604 218136 156656 218142
rect 156604 218078 156656 218084
rect 155224 213988 155276 213994
rect 155224 213930 155276 213936
rect 151176 149116 151228 149122
rect 151176 149058 151228 149064
rect 151084 128308 151136 128314
rect 151084 128250 151136 128256
rect 151084 125656 151136 125662
rect 151084 125598 151136 125604
rect 149796 121372 149848 121378
rect 149796 121314 149848 121320
rect 149796 114572 149848 114578
rect 149796 114514 149848 114520
rect 149704 77240 149756 77246
rect 149704 77182 149756 77188
rect 149808 73030 149836 114514
rect 151096 78674 151124 125598
rect 151188 90982 151216 149058
rect 151268 144968 151320 144974
rect 151268 144910 151320 144916
rect 151176 90976 151228 90982
rect 151176 90918 151228 90924
rect 151280 88262 151308 144910
rect 152464 143676 152516 143682
rect 152464 143618 152516 143624
rect 151360 128444 151412 128450
rect 151360 128386 151412 128392
rect 151268 88256 151320 88262
rect 151268 88198 151320 88204
rect 151372 80034 151400 128386
rect 152476 88330 152504 143618
rect 152556 139460 152608 139466
rect 152556 139402 152608 139408
rect 152464 88324 152516 88330
rect 152464 88266 152516 88272
rect 152568 85542 152596 139402
rect 152648 135380 152700 135386
rect 152648 135322 152700 135328
rect 152556 85536 152608 85542
rect 152556 85478 152608 85484
rect 152660 84182 152688 135322
rect 152740 132524 152792 132530
rect 152740 132466 152792 132472
rect 152648 84176 152700 84182
rect 152648 84118 152700 84124
rect 152752 82754 152780 132466
rect 155236 122806 155264 213930
rect 155316 164280 155368 164286
rect 155316 164222 155368 164228
rect 155224 122800 155276 122806
rect 155224 122742 155276 122748
rect 155328 97918 155356 164222
rect 155408 150476 155460 150482
rect 155408 150418 155460 150424
rect 155316 97912 155368 97918
rect 155316 97854 155368 97860
rect 155420 91050 155448 150418
rect 155500 146328 155552 146334
rect 155500 146270 155552 146276
rect 155408 91044 155460 91050
rect 155408 90986 155460 90992
rect 155512 89690 155540 146270
rect 156616 125594 156644 218078
rect 156696 189100 156748 189106
rect 156696 189042 156748 189048
rect 156604 125588 156656 125594
rect 156604 125530 156656 125536
rect 156708 110362 156736 189042
rect 156880 182232 156932 182238
rect 156880 182174 156932 182180
rect 156788 180940 156840 180946
rect 156788 180882 156840 180888
rect 156696 110356 156748 110362
rect 156696 110298 156748 110304
rect 156800 106282 156828 180882
rect 156892 107642 156920 182174
rect 156972 157480 157024 157486
rect 156972 157422 157024 157428
rect 156880 107636 156932 107642
rect 156880 107578 156932 107584
rect 156788 106276 156840 106282
rect 156788 106218 156840 106224
rect 156984 95198 157012 157422
rect 157996 129674 158024 225014
rect 162124 220856 162176 220862
rect 162124 220798 162176 220804
rect 160744 209908 160796 209914
rect 160744 209850 160796 209856
rect 159364 207052 159416 207058
rect 159364 206994 159416 207000
rect 158076 205692 158128 205698
rect 158076 205634 158128 205640
rect 157984 129668 158036 129674
rect 157984 129610 158036 129616
rect 158088 118658 158116 205634
rect 158168 168428 158220 168434
rect 158168 168370 158220 168376
rect 158076 118652 158128 118658
rect 158076 118594 158128 118600
rect 158180 100706 158208 168370
rect 158260 165640 158312 165646
rect 158260 165582 158312 165588
rect 158168 100700 158220 100706
rect 158168 100642 158220 100648
rect 158272 99278 158300 165582
rect 158352 160132 158404 160138
rect 158352 160074 158404 160080
rect 158260 99272 158312 99278
rect 158260 99214 158312 99220
rect 158364 96626 158392 160074
rect 159376 120018 159404 206994
rect 159456 197396 159508 197402
rect 159456 197338 159508 197344
rect 159364 120012 159416 120018
rect 159364 119954 159416 119960
rect 159468 114442 159496 197338
rect 159548 187808 159600 187814
rect 159548 187750 159600 187756
rect 159456 114436 159508 114442
rect 159456 114378 159508 114384
rect 159560 110294 159588 187750
rect 159640 165708 159692 165714
rect 159640 165650 159692 165656
rect 159548 110288 159600 110294
rect 159548 110230 159600 110236
rect 159652 100026 159680 165650
rect 160756 121446 160784 209850
rect 160836 172644 160888 172650
rect 160836 172586 160888 172592
rect 160744 121440 160796 121446
rect 160744 121382 160796 121388
rect 160848 102134 160876 172586
rect 160928 162920 160980 162926
rect 160928 162862 160980 162868
rect 160836 102128 160888 102134
rect 160836 102070 160888 102076
rect 159640 100020 159692 100026
rect 159640 99962 159692 99968
rect 160940 97986 160968 162862
rect 162136 126954 162164 220798
rect 166264 191276 166316 191282
rect 166264 191218 166316 191224
rect 164976 173936 165028 173942
rect 164976 173878 165028 173884
rect 162216 167068 162268 167074
rect 162216 167010 162268 167016
rect 162124 126948 162176 126954
rect 162124 126890 162176 126896
rect 162228 99346 162256 167010
rect 164884 133340 164936 133346
rect 164884 133282 164936 133288
rect 162216 99340 162268 99346
rect 162216 99282 162268 99288
rect 160928 97980 160980 97986
rect 160928 97922 160980 97928
rect 158352 96620 158404 96626
rect 158352 96562 158404 96568
rect 156972 95192 157024 95198
rect 156972 95134 157024 95140
rect 155500 89684 155552 89690
rect 155500 89626 155552 89632
rect 152740 82748 152792 82754
rect 152740 82690 152792 82696
rect 151360 80028 151412 80034
rect 151360 79970 151412 79976
rect 151084 78668 151136 78674
rect 151084 78610 151136 78616
rect 159364 75268 159416 75274
rect 159364 75210 159416 75216
rect 149796 73024 149848 73030
rect 149796 72966 149848 72972
rect 147128 69012 147180 69018
rect 147128 68954 147180 68960
rect 159376 62014 159404 75210
rect 159364 62008 159416 62014
rect 159364 61950 159416 61956
rect 146944 51060 146996 51066
rect 146944 51002 146996 51008
rect 144276 49632 144328 49638
rect 144276 49574 144328 49580
rect 142804 46912 142856 46918
rect 142804 46854 142856 46860
rect 141424 45484 141476 45490
rect 141424 45426 141476 45432
rect 140044 44056 140096 44062
rect 140044 43998 140096 44004
rect 133420 41336 133472 41342
rect 133420 41278 133472 41284
rect 164896 28558 164924 133282
rect 164988 103494 165016 173878
rect 164976 103488 165028 103494
rect 164976 103430 165028 103436
rect 166276 28694 166304 191218
rect 166356 150544 166408 150550
rect 166356 150486 166408 150492
rect 166368 92478 166396 150486
rect 169036 129742 169064 227734
rect 186318 227352 186374 227361
rect 186318 227287 186374 227296
rect 186332 226370 186360 227287
rect 186320 226364 186372 226370
rect 186320 226306 186372 226312
rect 186410 226264 186466 226273
rect 186410 226199 186466 226208
rect 186424 225078 186452 226199
rect 186412 225072 186464 225078
rect 186318 225040 186374 225049
rect 186412 225014 186464 225020
rect 186318 224975 186320 224984
rect 186372 224975 186374 224984
rect 186320 224946 186372 224952
rect 186318 223952 186374 223961
rect 186318 223887 186374 223896
rect 186332 223650 186360 223887
rect 186320 223644 186372 223650
rect 186320 223586 186372 223592
rect 186318 222728 186374 222737
rect 186318 222663 186374 222672
rect 186332 222222 186360 222663
rect 186320 222216 186372 222222
rect 186320 222158 186372 222164
rect 186318 221504 186374 221513
rect 186318 221439 186374 221448
rect 186332 220862 186360 221439
rect 186320 220856 186372 220862
rect 186320 220798 186372 220804
rect 186318 220416 186374 220425
rect 186318 220351 186374 220360
rect 186332 219502 186360 220351
rect 186320 219496 186372 219502
rect 186320 219438 186372 219444
rect 186410 219192 186466 219201
rect 186410 219127 186466 219136
rect 186424 218142 186452 219127
rect 186412 218136 186464 218142
rect 186318 218104 186374 218113
rect 186412 218078 186464 218084
rect 186318 218039 186320 218048
rect 186372 218039 186374 218048
rect 186320 218010 186372 218016
rect 186318 216880 186374 216889
rect 186318 216815 186374 216824
rect 186332 216714 186360 216815
rect 186320 216708 186372 216714
rect 186320 216650 186372 216656
rect 186318 215792 186374 215801
rect 186318 215727 186374 215736
rect 186332 215354 186360 215727
rect 186320 215348 186372 215354
rect 186320 215290 186372 215296
rect 186318 214568 186374 214577
rect 186318 214503 186374 214512
rect 186332 213994 186360 214503
rect 186320 213988 186372 213994
rect 186320 213930 186372 213936
rect 186318 213480 186374 213489
rect 186318 213415 186374 213424
rect 186332 212566 186360 213415
rect 186320 212560 186372 212566
rect 186320 212502 186372 212508
rect 186318 212256 186374 212265
rect 186318 212191 186374 212200
rect 186332 211206 186360 212191
rect 186320 211200 186372 211206
rect 186320 211142 186372 211148
rect 186410 211032 186466 211041
rect 186410 210967 186466 210976
rect 186318 209944 186374 209953
rect 186318 209879 186320 209888
rect 186372 209879 186374 209888
rect 186320 209850 186372 209856
rect 186424 209846 186452 210967
rect 186412 209840 186464 209846
rect 186412 209782 186464 209788
rect 186962 208720 187018 208729
rect 186962 208655 187018 208664
rect 186318 207632 186374 207641
rect 186318 207567 186374 207576
rect 186332 207058 186360 207567
rect 186320 207052 186372 207058
rect 186320 206994 186372 207000
rect 186318 206408 186374 206417
rect 186318 206343 186374 206352
rect 186332 205698 186360 206343
rect 186320 205692 186372 205698
rect 186320 205634 186372 205640
rect 186318 205320 186374 205329
rect 186318 205255 186374 205264
rect 186332 204338 186360 205255
rect 186320 204332 186372 204338
rect 186320 204274 186372 204280
rect 186410 204096 186466 204105
rect 186410 204031 186466 204040
rect 186318 203008 186374 203017
rect 186318 202943 186320 202952
rect 186372 202943 186374 202952
rect 186320 202914 186372 202920
rect 186424 202910 186452 204031
rect 186412 202904 186464 202910
rect 186412 202846 186464 202852
rect 186318 201784 186374 201793
rect 186318 201719 186374 201728
rect 186332 201550 186360 201719
rect 186320 201544 186372 201550
rect 186320 201486 186372 201492
rect 186318 200560 186374 200569
rect 186318 200495 186374 200504
rect 186332 200190 186360 200495
rect 186320 200184 186372 200190
rect 186320 200126 186372 200132
rect 186318 199472 186374 199481
rect 186318 199407 186374 199416
rect 186332 198762 186360 199407
rect 186320 198756 186372 198762
rect 186320 198698 186372 198704
rect 186318 198248 186374 198257
rect 186318 198183 186374 198192
rect 186332 197402 186360 198183
rect 186320 197396 186372 197402
rect 186320 197338 186372 197344
rect 186410 195936 186466 195945
rect 186410 195871 186466 195880
rect 186318 194848 186374 194857
rect 186318 194783 186374 194792
rect 186332 194682 186360 194783
rect 186320 194676 186372 194682
rect 186320 194618 186372 194624
rect 186424 194614 186452 195871
rect 186412 194608 186464 194614
rect 186412 194550 186464 194556
rect 186318 193624 186374 193633
rect 186318 193559 186374 193568
rect 186332 193254 186360 193559
rect 186320 193248 186372 193254
rect 186320 193190 186372 193196
rect 186318 192400 186374 192409
rect 186318 192335 186374 192344
rect 186332 191894 186360 192335
rect 186320 191888 186372 191894
rect 186320 191830 186372 191836
rect 186318 191312 186374 191321
rect 186318 191247 186374 191256
rect 186332 190534 186360 191247
rect 186320 190528 186372 190534
rect 186320 190470 186372 190476
rect 186318 190088 186374 190097
rect 186318 190023 186374 190032
rect 186332 189106 186360 190023
rect 186320 189100 186372 189106
rect 186320 189042 186372 189048
rect 186410 189000 186466 189009
rect 186410 188935 186466 188944
rect 186424 187814 186452 188935
rect 186412 187808 186464 187814
rect 186318 187776 186374 187785
rect 186412 187750 186464 187756
rect 186318 187711 186320 187720
rect 186372 187711 186374 187720
rect 186320 187682 186372 187688
rect 186318 186688 186374 186697
rect 186318 186623 186374 186632
rect 186332 186386 186360 186623
rect 186320 186380 186372 186386
rect 186320 186322 186372 186328
rect 186318 185464 186374 185473
rect 186318 185399 186374 185408
rect 186332 184958 186360 185399
rect 186320 184952 186372 184958
rect 186320 184894 186372 184900
rect 186318 184376 186374 184385
rect 186318 184311 186374 184320
rect 186332 183598 186360 184311
rect 186320 183592 186372 183598
rect 186320 183534 186372 183540
rect 186318 183152 186374 183161
rect 186318 183087 186374 183096
rect 186332 182238 186360 183087
rect 186320 182232 186372 182238
rect 186320 182174 186372 182180
rect 186410 181928 186466 181937
rect 186410 181863 186466 181872
rect 186320 180940 186372 180946
rect 186320 180882 186372 180888
rect 186332 180849 186360 180882
rect 186424 180878 186452 181863
rect 186412 180872 186464 180878
rect 186318 180840 186374 180849
rect 186412 180814 186464 180820
rect 186318 180775 186374 180784
rect 186318 179616 186374 179625
rect 186318 179551 186374 179560
rect 186332 179450 186360 179551
rect 186320 179444 186372 179450
rect 186320 179386 186372 179392
rect 186318 178528 186374 178537
rect 186318 178463 186374 178472
rect 186332 178090 186360 178463
rect 186320 178084 186372 178090
rect 186320 178026 186372 178032
rect 186318 177304 186374 177313
rect 186318 177239 186374 177248
rect 186332 176730 186360 177239
rect 186320 176724 186372 176730
rect 186320 176666 186372 176672
rect 186318 176216 186374 176225
rect 186318 176151 186374 176160
rect 186332 175302 186360 176151
rect 186320 175296 186372 175302
rect 186320 175238 186372 175244
rect 186318 174992 186374 175001
rect 186318 174927 186374 174936
rect 186332 173942 186360 174927
rect 186320 173936 186372 173942
rect 186320 173878 186372 173884
rect 186410 173768 186466 173777
rect 186410 173703 186466 173712
rect 186318 172680 186374 172689
rect 186318 172615 186320 172624
rect 186372 172615 186374 172624
rect 186320 172586 186372 172592
rect 186424 172582 186452 173703
rect 186412 172576 186464 172582
rect 186412 172518 186464 172524
rect 186318 171456 186374 171465
rect 186318 171391 186374 171400
rect 186332 171154 186360 171391
rect 186320 171148 186372 171154
rect 186320 171090 186372 171096
rect 186318 170368 186374 170377
rect 186318 170303 186374 170312
rect 186332 169794 186360 170303
rect 186320 169788 186372 169794
rect 186320 169730 186372 169736
rect 186318 169144 186374 169153
rect 186318 169079 186374 169088
rect 186332 168434 186360 169079
rect 186320 168428 186372 168434
rect 186320 168370 186372 168376
rect 186318 168056 186374 168065
rect 186318 167991 186374 168000
rect 186332 167074 186360 167991
rect 186320 167068 186372 167074
rect 186320 167010 186372 167016
rect 186410 166832 186466 166841
rect 186410 166767 186466 166776
rect 186318 165744 186374 165753
rect 186318 165679 186320 165688
rect 186372 165679 186374 165688
rect 186320 165650 186372 165656
rect 186424 165646 186452 166767
rect 186412 165640 186464 165646
rect 186412 165582 186464 165588
rect 186318 164520 186374 164529
rect 186318 164455 186374 164464
rect 186332 164286 186360 164455
rect 186320 164280 186372 164286
rect 186320 164222 186372 164228
rect 186318 163296 186374 163305
rect 186318 163231 186374 163240
rect 186332 162926 186360 163231
rect 186320 162920 186372 162926
rect 186320 162862 186372 162868
rect 186318 162208 186374 162217
rect 186318 162143 186374 162152
rect 186332 161498 186360 162143
rect 186320 161492 186372 161498
rect 186320 161434 186372 161440
rect 186318 160984 186374 160993
rect 186318 160919 186374 160928
rect 186332 160138 186360 160919
rect 186320 160132 186372 160138
rect 186320 160074 186372 160080
rect 186318 159896 186374 159905
rect 186318 159831 186374 159840
rect 186332 158778 186360 159831
rect 186320 158772 186372 158778
rect 186320 158714 186372 158720
rect 186410 158672 186466 158681
rect 186410 158607 186466 158616
rect 186318 157584 186374 157593
rect 186318 157519 186374 157528
rect 186332 157418 186360 157519
rect 186424 157486 186452 158607
rect 186412 157480 186464 157486
rect 186412 157422 186464 157428
rect 186320 157412 186372 157418
rect 186320 157354 186372 157360
rect 186318 156360 186374 156369
rect 186318 156295 186374 156304
rect 186332 155990 186360 156295
rect 186320 155984 186372 155990
rect 186320 155926 186372 155932
rect 186318 155272 186374 155281
rect 186318 155207 186374 155216
rect 186332 154630 186360 155207
rect 186320 154624 186372 154630
rect 186320 154566 186372 154572
rect 186318 154048 186374 154057
rect 186318 153983 186374 153992
rect 186332 153270 186360 153983
rect 186320 153264 186372 153270
rect 186320 153206 186372 153212
rect 186318 152824 186374 152833
rect 186318 152759 186374 152768
rect 186332 151842 186360 152759
rect 186320 151836 186372 151842
rect 186320 151778 186372 151784
rect 186410 151736 186466 151745
rect 186410 151671 186466 151680
rect 186424 150550 186452 151671
rect 186412 150544 186464 150550
rect 186318 150512 186374 150521
rect 186412 150486 186464 150492
rect 186318 150447 186320 150456
rect 186372 150447 186374 150456
rect 186320 150418 186372 150424
rect 186318 149424 186374 149433
rect 186318 149359 186374 149368
rect 186332 149122 186360 149359
rect 186320 149116 186372 149122
rect 186320 149058 186372 149064
rect 186318 148200 186374 148209
rect 186318 148135 186374 148144
rect 186332 147694 186360 148135
rect 186320 147688 186372 147694
rect 186320 147630 186372 147636
rect 186318 147112 186374 147121
rect 186318 147047 186374 147056
rect 186332 146334 186360 147047
rect 186320 146328 186372 146334
rect 186320 146270 186372 146276
rect 186318 145888 186374 145897
rect 186318 145823 186374 145832
rect 186332 144974 186360 145823
rect 186320 144968 186372 144974
rect 186320 144910 186372 144916
rect 186410 144664 186466 144673
rect 186410 144599 186466 144608
rect 186320 143676 186372 143682
rect 186320 143618 186372 143624
rect 186332 143585 186360 143618
rect 186424 143614 186452 144599
rect 186412 143608 186464 143614
rect 186318 143576 186374 143585
rect 186412 143550 186464 143556
rect 186318 143511 186374 143520
rect 186318 142352 186374 142361
rect 186318 142287 186374 142296
rect 186332 142186 186360 142287
rect 186320 142180 186372 142186
rect 186320 142122 186372 142128
rect 186318 140040 186374 140049
rect 186318 139975 186374 139984
rect 186332 139466 186360 139975
rect 186320 139460 186372 139466
rect 186320 139402 186372 139408
rect 186318 138952 186374 138961
rect 186318 138887 186374 138896
rect 186332 138038 186360 138887
rect 186320 138032 186372 138038
rect 186320 137974 186372 137980
rect 186318 137728 186374 137737
rect 186318 137663 186374 137672
rect 186332 136678 186360 137663
rect 186320 136672 186372 136678
rect 186320 136614 186372 136620
rect 186410 136640 186466 136649
rect 186410 136575 186466 136584
rect 186318 135416 186374 135425
rect 186424 135386 186452 136575
rect 186318 135351 186374 135360
rect 186412 135380 186464 135386
rect 186332 135318 186360 135351
rect 186412 135322 186464 135328
rect 186320 135312 186372 135318
rect 186320 135254 186372 135260
rect 186318 133104 186374 133113
rect 186318 133039 186374 133048
rect 186332 132530 186360 133039
rect 186320 132524 186372 132530
rect 186320 132466 186372 132472
rect 186318 131880 186374 131889
rect 186318 131815 186374 131824
rect 186332 131170 186360 131815
rect 186320 131164 186372 131170
rect 186320 131106 186372 131112
rect 186318 130792 186374 130801
rect 186318 130727 186374 130736
rect 186332 129810 186360 130727
rect 186320 129804 186372 129810
rect 186320 129746 186372 129752
rect 169024 129736 169076 129742
rect 169024 129678 169076 129684
rect 186410 129568 186466 129577
rect 186410 129503 186466 129512
rect 186318 128480 186374 128489
rect 186424 128450 186452 129503
rect 186318 128415 186374 128424
rect 186412 128444 186464 128450
rect 186332 128382 186360 128415
rect 186412 128386 186464 128392
rect 186320 128376 186372 128382
rect 186320 128318 186372 128324
rect 186318 127256 186374 127265
rect 186318 127191 186374 127200
rect 186332 127022 186360 127191
rect 186320 127016 186372 127022
rect 186320 126958 186372 126964
rect 186318 126032 186374 126041
rect 186318 125967 186374 125976
rect 186332 125662 186360 125967
rect 186320 125656 186372 125662
rect 186320 125598 186372 125604
rect 186318 124944 186374 124953
rect 186318 124879 186374 124888
rect 186332 124234 186360 124879
rect 186320 124228 186372 124234
rect 186320 124170 186372 124176
rect 186318 122632 186374 122641
rect 186318 122567 186374 122576
rect 186332 121514 186360 122567
rect 186320 121508 186372 121514
rect 186320 121450 186372 121456
rect 186410 121408 186466 121417
rect 186410 121343 186466 121352
rect 186318 120320 186374 120329
rect 186318 120255 186374 120264
rect 186332 120154 186360 120255
rect 186424 120222 186452 121343
rect 186412 120216 186464 120222
rect 186412 120158 186464 120164
rect 186320 120148 186372 120154
rect 186320 120090 186372 120096
rect 186976 120086 187004 208655
rect 409340 205601 409368 229066
rect 409892 209545 409920 279414
rect 409984 217297 410012 287642
rect 410064 282192 410116 282198
rect 410064 282134 410116 282140
rect 409970 217288 410026 217297
rect 409970 217223 410026 217232
rect 410076 213625 410104 282134
rect 411904 262948 411956 262954
rect 411904 262890 411956 262896
rect 411536 262880 411588 262886
rect 411536 262822 411588 262828
rect 410248 258800 410300 258806
rect 410248 258742 410300 258748
rect 410156 254652 410208 254658
rect 410156 254594 410208 254600
rect 410168 224369 410196 254594
rect 410260 228177 410288 258742
rect 411352 258732 411404 258738
rect 411352 258674 411404 258680
rect 410432 256080 410484 256086
rect 410432 256022 410484 256028
rect 410340 254720 410392 254726
rect 410340 254662 410392 254668
rect 410246 228168 410302 228177
rect 410246 228103 410302 228112
rect 410352 226273 410380 254662
rect 410444 231985 410472 256022
rect 411260 254584 411312 254590
rect 411260 254526 411312 254532
rect 410524 250640 410576 250646
rect 410524 250582 410576 250588
rect 410536 239601 410564 250582
rect 410522 239592 410578 239601
rect 410522 239527 410578 239536
rect 410430 231976 410486 231985
rect 410430 231911 410486 231920
rect 410338 226264 410394 226273
rect 410338 226199 410394 226208
rect 410154 224360 410210 224369
rect 410154 224295 410210 224304
rect 410062 213616 410118 213625
rect 410062 213551 410118 213560
rect 409878 209536 409934 209545
rect 409878 209471 409934 209480
rect 411272 207369 411300 254526
rect 411364 214849 411392 258674
rect 411444 256012 411496 256018
rect 411444 255954 411496 255960
rect 411350 214840 411406 214849
rect 411350 214775 411406 214784
rect 411456 211177 411484 255954
rect 411548 220561 411576 262822
rect 411628 261520 411680 261526
rect 411628 261462 411680 261468
rect 411640 230081 411668 261462
rect 411812 250572 411864 250578
rect 411812 250514 411864 250520
rect 411720 250504 411772 250510
rect 411720 250446 411772 250452
rect 411626 230072 411682 230081
rect 411626 230007 411682 230016
rect 411534 220552 411590 220561
rect 411534 220487 411590 220496
rect 411732 218657 411760 250446
rect 411824 222465 411852 250514
rect 411916 235793 411944 262890
rect 411902 235784 411958 235793
rect 411902 235719 411958 235728
rect 411810 222456 411866 222465
rect 411810 222391 411866 222400
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 411718 218648 411774 218657
rect 411718 218583 411774 218592
rect 580184 218074 580212 218991
rect 543004 218068 543056 218074
rect 543004 218010 543056 218016
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 411442 211168 411498 211177
rect 411442 211103 411498 211112
rect 411258 207360 411314 207369
rect 411258 207295 411314 207304
rect 409326 205592 409382 205601
rect 409326 205527 409382 205536
rect 411258 203552 411314 203561
rect 411258 203487 411314 203496
rect 411272 202910 411300 203487
rect 411260 202904 411312 202910
rect 411260 202846 411312 202852
rect 540244 202904 540296 202910
rect 540244 202846 540296 202852
rect 411258 201648 411314 201657
rect 411258 201583 411260 201592
rect 411312 201583 411314 201592
rect 414664 201612 414716 201618
rect 411260 201554 411312 201560
rect 414664 201554 414716 201560
rect 411258 199744 411314 199753
rect 411258 199679 411314 199688
rect 411272 198762 411300 199679
rect 411260 198756 411312 198762
rect 411260 198698 411312 198704
rect 411258 197840 411314 197849
rect 411258 197775 411314 197784
rect 411272 197402 411300 197775
rect 411260 197396 411312 197402
rect 411260 197338 411312 197344
rect 187054 197160 187110 197169
rect 187054 197095 187110 197104
rect 186964 120080 187016 120086
rect 186964 120022 187016 120028
rect 186318 119096 186374 119105
rect 186318 119031 186374 119040
rect 186332 118726 186360 119031
rect 186320 118720 186372 118726
rect 186320 118662 186372 118668
rect 186318 118008 186374 118017
rect 186318 117943 186374 117952
rect 186332 117366 186360 117943
rect 186320 117360 186372 117366
rect 186320 117302 186372 117308
rect 186318 116784 186374 116793
rect 186318 116719 186374 116728
rect 186332 116006 186360 116719
rect 186320 116000 186372 116006
rect 186320 115942 186372 115948
rect 186318 115560 186374 115569
rect 186318 115495 186374 115504
rect 186332 114578 186360 115495
rect 186320 114572 186372 114578
rect 186320 114514 186372 114520
rect 187068 114510 187096 197095
rect 411994 195936 412050 195945
rect 411994 195871 412050 195880
rect 411258 194032 411314 194041
rect 411258 193967 411314 193976
rect 411272 193594 411300 193967
rect 411260 193588 411312 193594
rect 411260 193530 411312 193536
rect 411902 192128 411958 192137
rect 411902 192063 411958 192072
rect 188344 191208 188396 191214
rect 188344 191150 188396 191156
rect 187146 141264 187202 141273
rect 187146 141199 187202 141208
rect 187056 114504 187108 114510
rect 187056 114446 187108 114452
rect 186962 113248 187018 113257
rect 186962 113183 187018 113192
rect 186318 112160 186374 112169
rect 186318 112095 186374 112104
rect 186332 111858 186360 112095
rect 186320 111852 186372 111858
rect 186320 111794 186372 111800
rect 186318 110936 186374 110945
rect 186318 110871 186374 110880
rect 186332 110498 186360 110871
rect 186320 110492 186372 110498
rect 186320 110434 186372 110440
rect 186318 109848 186374 109857
rect 186318 109783 186374 109792
rect 186332 109070 186360 109783
rect 186320 109064 186372 109070
rect 186320 109006 186372 109012
rect 186318 108624 186374 108633
rect 186318 108559 186374 108568
rect 186332 107710 186360 108559
rect 186320 107704 186372 107710
rect 186320 107646 186372 107652
rect 186410 107536 186466 107545
rect 186410 107471 186466 107480
rect 186424 106418 186452 107471
rect 186412 106412 186464 106418
rect 186412 106354 186464 106360
rect 186320 106344 186372 106350
rect 186318 106312 186320 106321
rect 186372 106312 186374 106321
rect 186318 106247 186374 106256
rect 186318 105088 186374 105097
rect 186318 105023 186374 105032
rect 186332 104922 186360 105023
rect 186320 104916 186372 104922
rect 186320 104858 186372 104864
rect 186318 104000 186374 104009
rect 186318 103935 186374 103944
rect 186332 103562 186360 103935
rect 186320 103556 186372 103562
rect 186320 103498 186372 103504
rect 186318 102776 186374 102785
rect 186318 102711 186374 102720
rect 186332 102202 186360 102711
rect 186320 102196 186372 102202
rect 186320 102138 186372 102144
rect 186318 101688 186374 101697
rect 186318 101623 186374 101632
rect 186332 100774 186360 101623
rect 186320 100768 186372 100774
rect 186320 100710 186372 100716
rect 186318 100464 186374 100473
rect 186318 100399 186374 100408
rect 186332 99414 186360 100399
rect 186320 99408 186372 99414
rect 186320 99350 186372 99356
rect 186410 99376 186466 99385
rect 186410 99311 186466 99320
rect 186318 98152 186374 98161
rect 186424 98122 186452 99311
rect 186318 98087 186374 98096
rect 186412 98116 186464 98122
rect 186332 98054 186360 98087
rect 186412 98058 186464 98064
rect 186320 98048 186372 98054
rect 186320 97990 186372 97996
rect 186318 96928 186374 96937
rect 186318 96863 186374 96872
rect 186332 96694 186360 96863
rect 186320 96688 186372 96694
rect 186320 96630 186372 96636
rect 186318 95840 186374 95849
rect 186318 95775 186374 95784
rect 186332 95266 186360 95775
rect 186320 95260 186372 95266
rect 186320 95202 186372 95208
rect 186318 94616 186374 94625
rect 186318 94551 186374 94560
rect 186332 93906 186360 94551
rect 186320 93900 186372 93906
rect 186320 93842 186372 93848
rect 186318 93528 186374 93537
rect 186318 93463 186374 93472
rect 186332 92546 186360 93463
rect 186320 92540 186372 92546
rect 186320 92482 186372 92488
rect 166356 92472 166408 92478
rect 166356 92414 166408 92420
rect 186318 91216 186374 91225
rect 186318 91151 186374 91160
rect 186332 91118 186360 91151
rect 181444 91112 181496 91118
rect 181444 91054 181496 91060
rect 186320 91112 186372 91118
rect 186320 91054 186372 91060
rect 181456 61946 181484 91054
rect 186318 89992 186374 90001
rect 186318 89927 186374 89936
rect 186332 89758 186360 89927
rect 186320 89752 186372 89758
rect 186320 89694 186372 89700
rect 186318 88904 186374 88913
rect 186318 88839 186374 88848
rect 186332 88398 186360 88839
rect 186320 88392 186372 88398
rect 186320 88334 186372 88340
rect 186318 87680 186374 87689
rect 186318 87615 186374 87624
rect 186332 87038 186360 87615
rect 186320 87032 186372 87038
rect 186320 86974 186372 86980
rect 186318 86456 186374 86465
rect 186318 86391 186374 86400
rect 186332 85610 186360 86391
rect 186320 85604 186372 85610
rect 186320 85546 186372 85552
rect 186410 84144 186466 84153
rect 186410 84079 186466 84088
rect 186318 83056 186374 83065
rect 186318 82991 186374 83000
rect 186332 82958 186360 82991
rect 186320 82952 186372 82958
rect 186320 82894 186372 82900
rect 186424 82890 186452 84079
rect 186412 82884 186464 82890
rect 186412 82826 186464 82832
rect 186318 80744 186374 80753
rect 186318 80679 186374 80688
rect 186332 80102 186360 80679
rect 186320 80096 186372 80102
rect 186320 80038 186372 80044
rect 186318 79520 186374 79529
rect 186318 79455 186374 79464
rect 186332 78742 186360 79455
rect 186320 78736 186372 78742
rect 186320 78678 186372 78684
rect 186410 77208 186466 77217
rect 186410 77143 186466 77152
rect 186320 76016 186372 76022
rect 186318 75984 186320 75993
rect 186372 75984 186374 75993
rect 186424 75954 186452 77143
rect 186318 75919 186374 75928
rect 186412 75948 186464 75954
rect 186412 75890 186464 75896
rect 186976 75206 187004 113183
rect 187160 86970 187188 141199
rect 187238 134192 187294 134201
rect 187238 134127 187294 134136
rect 187148 86964 187200 86970
rect 187148 86906 187200 86912
rect 187054 85368 187110 85377
rect 187054 85303 187110 85312
rect 186964 75200 187016 75206
rect 186964 75142 187016 75148
rect 186318 73672 186374 73681
rect 186318 73607 186374 73616
rect 186332 73234 186360 73607
rect 186320 73228 186372 73234
rect 186320 73170 186372 73176
rect 186318 72584 186374 72593
rect 186318 72519 186374 72528
rect 186332 71806 186360 72519
rect 181536 71800 181588 71806
rect 181536 71742 181588 71748
rect 186320 71800 186372 71806
rect 186320 71742 186372 71748
rect 181444 61940 181496 61946
rect 181444 61882 181496 61888
rect 181548 52426 181576 71742
rect 186318 71360 186374 71369
rect 186318 71295 186374 71304
rect 186332 70446 186360 71295
rect 186320 70440 186372 70446
rect 186320 70382 186372 70388
rect 186410 70272 186466 70281
rect 186410 70207 186466 70216
rect 186424 69154 186452 70207
rect 186412 69148 186464 69154
rect 186412 69090 186464 69096
rect 186320 69080 186372 69086
rect 186318 69048 186320 69057
rect 186372 69048 186374 69057
rect 186318 68983 186374 68992
rect 186318 67824 186374 67833
rect 186318 67759 186374 67768
rect 186332 67658 186360 67759
rect 181628 67652 181680 67658
rect 181628 67594 181680 67600
rect 186320 67652 186372 67658
rect 186320 67594 186372 67600
rect 181536 52420 181588 52426
rect 181536 52362 181588 52368
rect 181640 49706 181668 67594
rect 186318 66736 186374 66745
rect 186318 66671 186374 66680
rect 186332 66298 186360 66671
rect 186320 66292 186372 66298
rect 186320 66234 186372 66240
rect 186318 65512 186374 65521
rect 186318 65447 186374 65456
rect 186332 64938 186360 65447
rect 186320 64932 186372 64938
rect 186320 64874 186372 64880
rect 186318 64424 186374 64433
rect 186318 64359 186374 64368
rect 186332 63578 186360 64359
rect 181812 63572 181864 63578
rect 181812 63514 181864 63520
rect 186320 63572 186372 63578
rect 186320 63514 186372 63520
rect 181720 60852 181772 60858
rect 181720 60794 181772 60800
rect 181628 49700 181680 49706
rect 181628 49642 181680 49648
rect 181732 45422 181760 60794
rect 181824 48278 181852 63514
rect 186318 63200 186374 63209
rect 186318 63135 186374 63144
rect 186332 62150 186360 63135
rect 186320 62144 186372 62150
rect 186320 62086 186372 62092
rect 186410 62112 186466 62121
rect 186410 62047 186466 62056
rect 186318 60888 186374 60897
rect 186318 60823 186320 60832
rect 186372 60823 186374 60832
rect 186320 60794 186372 60800
rect 186424 60790 186452 62047
rect 186412 60784 186464 60790
rect 186412 60726 186464 60732
rect 186318 59800 186374 59809
rect 186318 59735 186374 59744
rect 186332 59430 186360 59735
rect 186320 59424 186372 59430
rect 186320 59366 186372 59372
rect 186318 58576 186374 58585
rect 186318 58511 186374 58520
rect 186332 58002 186360 58511
rect 186320 57996 186372 58002
rect 186320 57938 186372 57944
rect 187068 57934 187096 85303
rect 187252 82822 187280 134127
rect 187330 123720 187386 123729
rect 187330 123655 187386 123664
rect 187240 82816 187292 82822
rect 187240 82758 187292 82764
rect 187146 81832 187202 81841
rect 187146 81767 187202 81776
rect 187056 57928 187108 57934
rect 187056 57870 187108 57876
rect 186962 57352 187018 57361
rect 186962 57287 187018 57296
rect 186318 56264 186374 56273
rect 186318 56199 186374 56208
rect 186332 55282 186360 56199
rect 186320 55276 186372 55282
rect 186320 55218 186372 55224
rect 186318 55040 186374 55049
rect 186318 54975 186374 54984
rect 186332 53854 186360 54975
rect 186320 53848 186372 53854
rect 186320 53790 186372 53796
rect 186318 52728 186374 52737
rect 186318 52663 186374 52672
rect 186332 52494 186360 52663
rect 186320 52488 186372 52494
rect 186320 52430 186372 52436
rect 186318 51640 186374 51649
rect 186318 51575 186374 51584
rect 186332 51134 186360 51575
rect 186320 51128 186372 51134
rect 186320 51070 186372 51076
rect 186318 49192 186374 49201
rect 186318 49127 186374 49136
rect 186332 48346 186360 49127
rect 186320 48340 186372 48346
rect 186320 48282 186372 48288
rect 181812 48272 181864 48278
rect 181812 48214 181864 48220
rect 186318 48104 186374 48113
rect 186318 48039 186374 48048
rect 186332 46986 186360 48039
rect 186320 46980 186372 46986
rect 186320 46922 186372 46928
rect 181720 45416 181772 45422
rect 181720 45358 181772 45364
rect 186318 44568 186374 44577
rect 186318 44503 186374 44512
rect 186332 44198 186360 44503
rect 182088 44192 182140 44198
rect 182088 44134 182140 44140
rect 186320 44192 186372 44198
rect 186320 44134 186372 44140
rect 182100 39370 182128 44134
rect 186976 44130 187004 57287
rect 187160 56574 187188 81767
rect 187344 77994 187372 123655
rect 187422 114472 187478 114481
rect 187422 114407 187478 114416
rect 187436 101454 187464 114407
rect 187424 101448 187476 101454
rect 187424 101390 187476 101396
rect 187514 92304 187570 92313
rect 187514 92239 187570 92248
rect 187422 78296 187478 78305
rect 187422 78231 187478 78240
rect 187332 77988 187384 77994
rect 187332 77930 187384 77936
rect 187238 74896 187294 74905
rect 187238 74831 187294 74840
rect 187148 56568 187200 56574
rect 187148 56510 187200 56516
rect 187054 53952 187110 53961
rect 187054 53887 187110 53896
rect 186964 44124 187016 44130
rect 186964 44066 187016 44072
rect 186318 43480 186374 43489
rect 186318 43415 186374 43424
rect 186332 42838 186360 43415
rect 186320 42832 186372 42838
rect 186320 42774 186372 42780
rect 187068 42770 187096 53887
rect 187252 53786 187280 74831
rect 187436 55894 187464 78231
rect 187528 75274 187556 92239
rect 187516 75268 187568 75274
rect 187516 75210 187568 75216
rect 187424 55888 187476 55894
rect 187424 55830 187476 55836
rect 187240 53780 187292 53786
rect 187240 53722 187292 53728
rect 187146 50416 187202 50425
rect 187146 50351 187202 50360
rect 187056 42764 187108 42770
rect 187056 42706 187108 42712
rect 186410 42256 186466 42265
rect 186410 42191 186466 42200
rect 182088 39364 182140 39370
rect 182088 39306 182140 39312
rect 186318 38720 186374 38729
rect 186318 38655 186320 38664
rect 186372 38655 186374 38664
rect 186320 38626 186372 38632
rect 186318 37632 186374 37641
rect 186318 37567 186374 37576
rect 186332 37330 186360 37567
rect 186320 37324 186372 37330
rect 186320 37266 186372 37272
rect 186424 37262 186452 42191
rect 187160 41410 187188 50351
rect 187422 46880 187478 46889
rect 187422 46815 187478 46824
rect 187238 45792 187294 45801
rect 187238 45727 187294 45736
rect 187148 41404 187200 41410
rect 187148 41346 187200 41352
rect 186962 41168 187018 41177
rect 186962 41103 187018 41112
rect 186412 37256 186464 37262
rect 186412 37198 186464 37204
rect 186318 36408 186374 36417
rect 186318 36343 186374 36352
rect 186332 35970 186360 36343
rect 186320 35964 186372 35970
rect 186320 35906 186372 35912
rect 186976 35902 187004 41103
rect 187054 39944 187110 39953
rect 187054 39879 187110 39888
rect 186964 35896 187016 35902
rect 186964 35838 187016 35844
rect 187068 35834 187096 39879
rect 187252 38554 187280 45727
rect 187436 38622 187464 46815
rect 187424 38616 187476 38622
rect 187424 38558 187476 38564
rect 187240 38548 187292 38554
rect 187240 38490 187292 38496
rect 187056 35828 187108 35834
rect 187056 35770 187108 35776
rect 186410 35320 186466 35329
rect 186410 35255 186466 35264
rect 186318 34096 186374 34105
rect 186318 34031 186374 34040
rect 186332 33182 186360 34031
rect 186320 33176 186372 33182
rect 186320 33118 186372 33124
rect 186424 33114 186452 35255
rect 186412 33108 186464 33114
rect 186412 33050 186464 33056
rect 186410 33008 186466 33017
rect 186410 32943 186466 32952
rect 186424 31890 186452 32943
rect 186412 31884 186464 31890
rect 186412 31826 186464 31832
rect 186320 31816 186372 31822
rect 186318 31784 186320 31793
rect 186372 31784 186374 31793
rect 186318 31719 186374 31728
rect 186320 31068 186372 31074
rect 186320 31010 186372 31016
rect 186332 30705 186360 31010
rect 186318 30696 186374 30705
rect 186318 30631 186374 30640
rect 166264 28688 166316 28694
rect 166264 28630 166316 28636
rect 164884 28552 164936 28558
rect 164884 28494 164936 28500
rect 188356 28490 188384 191150
rect 189724 191140 189776 191146
rect 189724 191082 189776 191088
rect 188528 133272 188580 133278
rect 188528 133214 188580 133220
rect 188436 133204 188488 133210
rect 188436 133146 188488 133152
rect 188448 28762 188476 133146
rect 188540 28830 188568 133214
rect 188528 28824 188580 28830
rect 188528 28766 188580 28772
rect 188436 28756 188488 28762
rect 188436 28698 188488 28704
rect 188344 28484 188396 28490
rect 188344 28426 188396 28432
rect 133144 28348 133196 28354
rect 133144 28290 133196 28296
rect 189736 28218 189764 191082
rect 411258 190224 411314 190233
rect 411258 190159 411314 190168
rect 411272 189106 411300 190159
rect 411260 189100 411312 189106
rect 411260 189042 411312 189048
rect 411258 188320 411314 188329
rect 411258 188255 411314 188264
rect 411272 187746 411300 188255
rect 411260 187740 411312 187746
rect 411260 187682 411312 187688
rect 411258 186416 411314 186425
rect 411258 186351 411260 186360
rect 411312 186351 411314 186360
rect 411260 186322 411312 186328
rect 411258 184512 411314 184521
rect 411258 184447 411314 184456
rect 411272 183598 411300 184447
rect 411260 183592 411312 183598
rect 411260 183534 411312 183540
rect 411258 182608 411314 182617
rect 411258 182543 411314 182552
rect 411272 182238 411300 182543
rect 411260 182232 411312 182238
rect 411260 182174 411312 182180
rect 411258 180704 411314 180713
rect 411258 180639 411314 180648
rect 411272 179450 411300 180639
rect 411260 179444 411312 179450
rect 411260 179386 411312 179392
rect 411258 178800 411314 178809
rect 411258 178735 411314 178744
rect 411272 178090 411300 178735
rect 411260 178084 411312 178090
rect 411260 178026 411312 178032
rect 411258 177032 411314 177041
rect 411258 176967 411314 176976
rect 411272 176730 411300 176967
rect 411260 176724 411312 176730
rect 411260 176666 411312 176672
rect 411258 175128 411314 175137
rect 411258 175063 411314 175072
rect 411272 174486 411300 175063
rect 411260 174480 411312 174486
rect 411260 174422 411312 174428
rect 411258 173224 411314 173233
rect 411258 173159 411314 173168
rect 411272 172582 411300 173159
rect 411260 172576 411312 172582
rect 411260 172518 411312 172524
rect 411258 171320 411314 171329
rect 411258 171255 411314 171264
rect 411272 171154 411300 171255
rect 411260 171148 411312 171154
rect 411260 171090 411312 171096
rect 411258 169416 411314 169425
rect 411258 169351 411314 169360
rect 411272 168434 411300 169351
rect 411260 168428 411312 168434
rect 411260 168370 411312 168376
rect 411258 167512 411314 167521
rect 411258 167447 411314 167456
rect 411272 167074 411300 167447
rect 411260 167068 411312 167074
rect 411260 167010 411312 167016
rect 411258 165608 411314 165617
rect 411258 165543 411314 165552
rect 411272 164286 411300 165543
rect 411260 164280 411312 164286
rect 411260 164222 411312 164228
rect 411258 163704 411314 163713
rect 411258 163639 411314 163648
rect 411272 162926 411300 163639
rect 411260 162920 411312 162926
rect 411260 162862 411312 162868
rect 411258 161800 411314 161809
rect 411258 161735 411314 161744
rect 411272 161498 411300 161735
rect 411260 161492 411312 161498
rect 411260 161434 411312 161440
rect 411258 159896 411314 159905
rect 411258 159831 411314 159840
rect 411272 158778 411300 159831
rect 411260 158772 411312 158778
rect 411260 158714 411312 158720
rect 411258 157992 411314 158001
rect 411258 157927 411314 157936
rect 411272 157418 411300 157927
rect 411260 157412 411312 157418
rect 411260 157354 411312 157360
rect 411258 156088 411314 156097
rect 411258 156023 411314 156032
rect 411272 155990 411300 156023
rect 411260 155984 411312 155990
rect 411260 155926 411312 155932
rect 411258 154184 411314 154193
rect 411258 154119 411314 154128
rect 411272 153270 411300 154119
rect 411260 153264 411312 153270
rect 411260 153206 411312 153212
rect 411258 152280 411314 152289
rect 411258 152215 411314 152224
rect 411272 151842 411300 152215
rect 411260 151836 411312 151842
rect 411260 151778 411312 151784
rect 411258 150376 411314 150385
rect 411258 150311 411314 150320
rect 411272 149122 411300 150311
rect 411260 149116 411312 149122
rect 411260 149058 411312 149064
rect 411258 148472 411314 148481
rect 411258 148407 411314 148416
rect 411272 147694 411300 148407
rect 411260 147688 411312 147694
rect 411260 147630 411312 147636
rect 411258 146568 411314 146577
rect 411258 146503 411314 146512
rect 411272 146334 411300 146503
rect 411260 146328 411312 146334
rect 411260 146270 411312 146276
rect 411258 144664 411314 144673
rect 411258 144599 411314 144608
rect 411272 143614 411300 144599
rect 411260 143608 411312 143614
rect 411260 143550 411312 143556
rect 411258 142760 411314 142769
rect 411258 142695 411314 142704
rect 411272 142186 411300 142695
rect 411260 142180 411312 142186
rect 411260 142122 411312 142128
rect 411258 140992 411314 141001
rect 411258 140927 411314 140936
rect 411272 140826 411300 140927
rect 411260 140820 411312 140826
rect 411260 140762 411312 140768
rect 411258 139088 411314 139097
rect 411258 139023 411314 139032
rect 411272 138038 411300 139023
rect 411260 138032 411312 138038
rect 411260 137974 411312 137980
rect 411258 137184 411314 137193
rect 411258 137119 411314 137128
rect 411272 136678 411300 137119
rect 411260 136672 411312 136678
rect 411260 136614 411312 136620
rect 411260 135312 411312 135318
rect 411258 135280 411260 135289
rect 411312 135280 411314 135289
rect 411258 135215 411314 135224
rect 411258 133376 411314 133385
rect 411258 133311 411314 133320
rect 411272 132530 411300 133311
rect 411260 132524 411312 132530
rect 411260 132466 411312 132472
rect 190000 131912 190052 131918
rect 190000 131854 190052 131860
rect 189908 131844 189960 131850
rect 189908 131786 189960 131792
rect 189816 131776 189868 131782
rect 189816 131718 189868 131724
rect 189724 28212 189776 28218
rect 189724 28154 189776 28160
rect 189828 28150 189856 131718
rect 189920 28422 189948 131786
rect 190012 28626 190040 131854
rect 411258 131472 411314 131481
rect 411258 131407 411314 131416
rect 411272 131170 411300 131407
rect 411260 131164 411312 131170
rect 411260 131106 411312 131112
rect 190184 130484 190236 130490
rect 190184 130426 190236 130432
rect 190092 130416 190144 130422
rect 190092 130358 190144 130364
rect 190000 28620 190052 28626
rect 190000 28562 190052 28568
rect 189908 28416 189960 28422
rect 189908 28358 189960 28364
rect 190104 28286 190132 130358
rect 190092 28280 190144 28286
rect 190092 28222 190144 28228
rect 189816 28144 189868 28150
rect 189816 28086 189868 28092
rect 190196 28082 190224 130426
rect 411258 129568 411314 129577
rect 411258 129503 411314 129512
rect 411272 128518 411300 129503
rect 411260 128512 411312 128518
rect 411260 128454 411312 128460
rect 411258 127664 411314 127673
rect 411258 127599 411314 127608
rect 411272 127090 411300 127599
rect 411260 127084 411312 127090
rect 411260 127026 411312 127032
rect 411258 125760 411314 125769
rect 411258 125695 411260 125704
rect 411312 125695 411314 125704
rect 411260 125666 411312 125672
rect 411258 123856 411314 123865
rect 411258 123791 411314 123800
rect 411272 122874 411300 123791
rect 411260 122868 411312 122874
rect 411260 122810 411312 122816
rect 411258 121952 411314 121961
rect 411258 121887 411314 121896
rect 411272 121582 411300 121887
rect 411260 121576 411312 121582
rect 411260 121518 411312 121524
rect 411258 120048 411314 120057
rect 411258 119983 411314 119992
rect 411272 118726 411300 119983
rect 411260 118720 411312 118726
rect 411260 118662 411312 118668
rect 411258 118144 411314 118153
rect 411258 118079 411314 118088
rect 411272 117366 411300 118079
rect 411260 117360 411312 117366
rect 411260 117302 411312 117308
rect 411258 116240 411314 116249
rect 411258 116175 411314 116184
rect 411272 116006 411300 116175
rect 411260 116000 411312 116006
rect 411260 115942 411312 115948
rect 411916 115938 411944 192063
rect 412008 120086 412036 195871
rect 413376 193588 413428 193594
rect 413376 193530 413428 193536
rect 412272 129804 412324 129810
rect 412272 129746 412324 129752
rect 411996 120080 412048 120086
rect 411996 120022 412048 120028
rect 411904 115932 411956 115938
rect 411904 115874 411956 115880
rect 411994 114336 412050 114345
rect 411994 114271 412050 114280
rect 411258 112432 411314 112441
rect 411258 112367 411314 112376
rect 411272 111858 411300 112367
rect 411260 111852 411312 111858
rect 411260 111794 411312 111800
rect 411258 110528 411314 110537
rect 411258 110463 411260 110472
rect 411312 110463 411314 110472
rect 411260 110434 411312 110440
rect 411902 108624 411958 108633
rect 411902 108559 411958 108568
rect 411258 106720 411314 106729
rect 411258 106655 411314 106664
rect 411272 106350 411300 106655
rect 411260 106344 411312 106350
rect 411260 106286 411312 106292
rect 411258 104816 411314 104825
rect 411258 104751 411314 104760
rect 411272 103562 411300 104751
rect 411260 103556 411312 103562
rect 411260 103498 411312 103504
rect 411258 103048 411314 103057
rect 411258 102983 411314 102992
rect 411272 102202 411300 102983
rect 411260 102196 411312 102202
rect 411260 102138 411312 102144
rect 411258 101144 411314 101153
rect 411258 101079 411314 101088
rect 411272 100774 411300 101079
rect 411260 100768 411312 100774
rect 411260 100710 411312 100716
rect 411258 99240 411314 99249
rect 411258 99175 411314 99184
rect 411272 98054 411300 99175
rect 411260 98048 411312 98054
rect 411260 97990 411312 97996
rect 411810 95432 411866 95441
rect 411810 95367 411866 95376
rect 411350 93528 411406 93537
rect 411350 93463 411406 93472
rect 411364 92546 411392 93463
rect 411352 92540 411404 92546
rect 411352 92482 411404 92488
rect 411260 92472 411312 92478
rect 411260 92414 411312 92420
rect 411272 91633 411300 92414
rect 411258 91624 411314 91633
rect 411258 91559 411314 91568
rect 410524 91044 410576 91050
rect 410524 90986 410576 90992
rect 195256 30110 195454 30138
rect 206296 30110 206402 30138
rect 217442 30110 217824 30138
rect 195256 28898 195284 30110
rect 206296 29170 206324 30110
rect 206284 29164 206336 29170
rect 206284 29106 206336 29112
rect 206296 29034 206324 29106
rect 217796 29034 217824 30110
rect 227732 30110 228390 30138
rect 239048 30110 239430 30138
rect 250088 30110 250378 30138
rect 261128 30110 261418 30138
rect 271984 30110 272366 30138
rect 283024 30110 283406 30138
rect 294064 30110 294354 30138
rect 316236 30110 316434 30138
rect 327092 30110 327382 30138
rect 338132 30110 338422 30138
rect 349172 30110 349370 30138
rect 360212 30110 360410 30138
rect 371252 30110 371358 30138
rect 382292 30110 382398 30138
rect 393346 30110 393452 30138
rect 404386 30110 404492 30138
rect 205640 29028 205692 29034
rect 205640 28970 205692 28976
rect 206284 29028 206336 29034
rect 206284 28970 206336 28976
rect 217784 29028 217836 29034
rect 217784 28970 217836 28976
rect 195244 28892 195296 28898
rect 195244 28834 195296 28840
rect 190184 28076 190236 28082
rect 190184 28018 190236 28024
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 1308 4072 1360 4078
rect 1308 4014 1360 4020
rect 1320 3670 1348 4014
rect 2700 3738 2728 4082
rect 195256 4078 195284 28834
rect 205652 4146 205680 28970
rect 227732 6866 227760 30110
rect 239048 28354 239076 30110
rect 239036 28348 239088 28354
rect 239036 28290 239088 28296
rect 250088 28082 250116 30110
rect 261128 28150 261156 30110
rect 271984 28218 272012 30110
rect 283024 29306 283052 30110
rect 283012 29300 283064 29306
rect 283012 29242 283064 29248
rect 294064 28286 294092 30110
rect 316236 29238 316264 30110
rect 316224 29232 316276 29238
rect 316224 29174 316276 29180
rect 327092 28422 327120 30110
rect 338132 28490 338160 30110
rect 349172 28558 349200 30110
rect 360212 28694 360240 30110
rect 371252 29102 371280 30110
rect 371240 29096 371292 29102
rect 371240 29038 371292 29044
rect 360200 28688 360252 28694
rect 360200 28630 360252 28636
rect 382292 28626 382320 30110
rect 393424 28762 393452 30110
rect 404464 28830 404492 30110
rect 410536 29170 410564 90986
rect 411258 89720 411314 89729
rect 411258 89655 411260 89664
rect 411312 89655 411314 89664
rect 411260 89626 411312 89632
rect 411824 89010 411852 95367
rect 411812 89004 411864 89010
rect 411812 88946 411864 88952
rect 411260 88324 411312 88330
rect 411260 88266 411312 88272
rect 411272 87825 411300 88266
rect 411258 87816 411314 87825
rect 411258 87751 411314 87760
rect 411260 86964 411312 86970
rect 411260 86906 411312 86912
rect 411272 85921 411300 86906
rect 411258 85912 411314 85921
rect 411258 85847 411314 85856
rect 411258 84008 411314 84017
rect 411258 83943 411314 83952
rect 411272 82890 411300 83943
rect 411260 82884 411312 82890
rect 411260 82826 411312 82832
rect 411258 80200 411314 80209
rect 411258 80135 411260 80144
rect 411312 80135 411314 80144
rect 411260 80106 411312 80112
rect 411260 78328 411312 78334
rect 411258 78296 411260 78305
rect 411312 78296 411314 78305
rect 411258 78231 411314 78240
rect 411260 77240 411312 77246
rect 411260 77182 411312 77188
rect 411272 76401 411300 77182
rect 411258 76392 411314 76401
rect 411258 76327 411314 76336
rect 411260 74520 411312 74526
rect 411258 74488 411260 74497
rect 411312 74488 411314 74497
rect 411258 74423 411314 74432
rect 411260 72820 411312 72826
rect 411260 72762 411312 72768
rect 411272 72593 411300 72762
rect 411258 72584 411314 72593
rect 411258 72519 411314 72528
rect 411350 68776 411406 68785
rect 411350 68711 411406 68720
rect 411364 67658 411392 68711
rect 411352 67652 411404 67658
rect 411352 67594 411404 67600
rect 411260 67584 411312 67590
rect 411260 67526 411312 67532
rect 411272 67017 411300 67526
rect 411258 67008 411314 67017
rect 411258 66943 411314 66952
rect 411258 65104 411314 65113
rect 411258 65039 411260 65048
rect 411312 65039 411314 65048
rect 411260 65010 411312 65016
rect 411260 63504 411312 63510
rect 411260 63446 411312 63452
rect 411272 63209 411300 63446
rect 411258 63200 411314 63209
rect 411258 63135 411314 63144
rect 411258 61296 411314 61305
rect 411258 61231 411314 61240
rect 411272 60790 411300 61231
rect 411260 60784 411312 60790
rect 411260 60726 411312 60732
rect 411352 60716 411404 60722
rect 411352 60658 411404 60664
rect 411364 59401 411392 60658
rect 411350 59392 411406 59401
rect 411350 59327 411406 59336
rect 411260 57860 411312 57866
rect 411260 57802 411312 57808
rect 411272 57497 411300 57802
rect 411258 57488 411314 57497
rect 411258 57423 411314 57432
rect 411258 55584 411314 55593
rect 411258 55519 411314 55528
rect 411272 55282 411300 55519
rect 411260 55276 411312 55282
rect 411260 55218 411312 55224
rect 411260 50992 411312 50998
rect 411260 50934 411312 50940
rect 411272 49881 411300 50934
rect 411258 49872 411314 49881
rect 411258 49807 411314 49816
rect 411260 48068 411312 48074
rect 411260 48010 411312 48016
rect 411272 47977 411300 48010
rect 411258 47968 411314 47977
rect 411258 47903 411314 47912
rect 411258 46064 411314 46073
rect 411258 45999 411314 46008
rect 411272 45626 411300 45999
rect 411260 45620 411312 45626
rect 411260 45562 411312 45568
rect 411810 44160 411866 44169
rect 411810 44095 411866 44104
rect 411260 42560 411312 42566
rect 411260 42502 411312 42508
rect 411272 42265 411300 42502
rect 411258 42256 411314 42265
rect 411258 42191 411314 42200
rect 411260 41404 411312 41410
rect 411260 41346 411312 41352
rect 411272 40361 411300 41346
rect 411258 40352 411314 40361
rect 411258 40287 411314 40296
rect 411260 38616 411312 38622
rect 411260 38558 411312 38564
rect 411272 38457 411300 38558
rect 411258 38448 411314 38457
rect 411258 38383 411314 38392
rect 411260 37256 411312 37262
rect 411260 37198 411312 37204
rect 411272 36553 411300 37198
rect 411258 36544 411314 36553
rect 411258 36479 411314 36488
rect 411260 35828 411312 35834
rect 411260 35770 411312 35776
rect 411272 34649 411300 35770
rect 411258 34640 411314 34649
rect 411258 34575 411314 34584
rect 411260 33040 411312 33046
rect 411260 32982 411312 32988
rect 411272 32745 411300 32982
rect 411258 32736 411314 32745
rect 411258 32671 411314 32680
rect 411824 31754 411852 44095
rect 411916 42770 411944 108559
rect 412008 48278 412036 114271
rect 412086 97336 412142 97345
rect 412086 97271 412142 97280
rect 411996 48272 412048 48278
rect 411996 48214 412048 48220
rect 411904 42764 411956 42770
rect 411904 42706 411956 42712
rect 412100 33114 412128 97271
rect 412180 89004 412232 89010
rect 412180 88946 412232 88952
rect 412088 33108 412140 33114
rect 412088 33050 412140 33056
rect 411812 31748 411864 31754
rect 411812 31690 411864 31696
rect 412192 31550 412220 88946
rect 412284 84194 412312 129746
rect 412364 128376 412416 128382
rect 412364 128318 412416 128324
rect 412376 93854 412404 128318
rect 413284 121508 413336 121514
rect 413284 121450 413336 121456
rect 412376 93826 412496 93854
rect 412284 84166 412404 84194
rect 412376 70689 412404 84166
rect 412468 82113 412496 93826
rect 412454 82104 412510 82113
rect 412454 82039 412510 82048
rect 412362 70680 412418 70689
rect 412362 70615 412418 70624
rect 412270 53680 412326 53689
rect 412270 53615 412326 53624
rect 412284 31686 412312 53615
rect 412362 51776 412418 51785
rect 412362 51711 412418 51720
rect 412272 31680 412324 31686
rect 412272 31622 412324 31628
rect 412376 31618 412404 51711
rect 413296 38622 413324 121450
rect 413388 118658 413416 193530
rect 414676 139398 414704 201554
rect 428464 189100 428516 189106
rect 428464 189042 428516 189048
rect 418988 186380 419040 186386
rect 418988 186322 419040 186328
rect 417424 176724 417476 176730
rect 417424 176666 417476 176672
rect 414940 174480 414992 174486
rect 414940 174422 414992 174428
rect 414664 139392 414716 139398
rect 414664 139334 414716 139340
rect 413468 131504 413520 131510
rect 413468 131446 413520 131452
rect 413376 118652 413428 118658
rect 413376 118594 413428 118600
rect 413376 103556 413428 103562
rect 413376 103498 413428 103504
rect 413388 40050 413416 103498
rect 413480 72826 413508 131446
rect 414664 131368 414716 131374
rect 414664 131310 414716 131316
rect 413560 127016 413612 127022
rect 413560 126958 413612 126964
rect 413572 89690 413600 126958
rect 413652 125656 413704 125662
rect 413652 125598 413704 125604
rect 413560 89684 413612 89690
rect 413560 89626 413612 89632
rect 413560 80164 413612 80170
rect 413560 80106 413612 80112
rect 413468 72820 413520 72826
rect 413468 72762 413520 72768
rect 413468 65068 413520 65074
rect 413468 65010 413520 65016
rect 413376 40044 413428 40050
rect 413376 39986 413428 39992
rect 413284 38616 413336 38622
rect 413284 38558 413336 38564
rect 412364 31612 412416 31618
rect 412364 31554 412416 31560
rect 412180 31544 412232 31550
rect 412180 31486 412232 31492
rect 411258 30968 411314 30977
rect 411258 30903 411314 30912
rect 410524 29164 410576 29170
rect 410524 29106 410576 29112
rect 404452 28824 404504 28830
rect 404452 28766 404504 28772
rect 393412 28756 393464 28762
rect 393412 28698 393464 28704
rect 411272 28694 411300 30903
rect 413480 28830 413508 65010
rect 413572 29102 413600 80106
rect 413664 78334 413692 125598
rect 414020 96076 414072 96082
rect 414020 96018 414072 96024
rect 414032 91118 414060 96018
rect 414020 91112 414072 91118
rect 414020 91054 414072 91060
rect 413652 78328 413704 78334
rect 413652 78270 413704 78276
rect 414676 42566 414704 131310
rect 414756 131300 414808 131306
rect 414756 131242 414808 131248
rect 414768 50998 414796 131242
rect 414848 124228 414900 124234
rect 414848 124170 414900 124176
rect 414756 50992 414808 50998
rect 414756 50934 414808 50940
rect 414860 48074 414888 124170
rect 414952 102134 414980 174422
rect 415032 131164 415084 131170
rect 415032 131106 415084 131112
rect 414940 102128 414992 102134
rect 414940 102070 414992 102076
rect 414940 98048 414992 98054
rect 414940 97990 414992 97996
rect 414848 48068 414900 48074
rect 414848 48010 414900 48016
rect 414664 42560 414716 42566
rect 414664 42502 414716 42508
rect 414952 34474 414980 97990
rect 415044 90370 415072 131106
rect 416044 125724 416096 125730
rect 416044 125666 416096 125672
rect 415952 99408 416004 99414
rect 415952 99350 416004 99356
rect 415964 96082 415992 99350
rect 415952 96076 416004 96082
rect 415952 96018 416004 96024
rect 415032 90364 415084 90370
rect 415032 90306 415084 90312
rect 416056 57934 416084 125666
rect 416136 121576 416188 121582
rect 416136 121518 416188 121524
rect 416044 57928 416096 57934
rect 416044 57870 416096 57876
rect 416148 55214 416176 121518
rect 417436 103494 417464 176666
rect 417516 153264 417568 153270
rect 417516 153206 417568 153212
rect 417424 103488 417476 103494
rect 417424 103430 417476 103436
rect 417424 100768 417476 100774
rect 417424 100710 417476 100716
rect 416136 55208 416188 55214
rect 416136 55150 416188 55156
rect 417436 35902 417464 100710
rect 417528 82822 417556 153206
rect 417608 149116 417660 149122
rect 417608 149058 417660 149064
rect 417516 82816 417568 82822
rect 417516 82758 417568 82764
rect 417620 80034 417648 149058
rect 417700 140820 417752 140826
rect 417700 140762 417752 140768
rect 417608 80028 417660 80034
rect 417608 79970 417660 79976
rect 417712 71738 417740 140762
rect 418804 129872 418856 129878
rect 418804 129814 418856 129820
rect 418160 106752 418212 106758
rect 418160 106694 418212 106700
rect 417792 106344 417844 106350
rect 417792 106286 417844 106292
rect 417700 71732 417752 71738
rect 417700 71674 417752 71680
rect 417804 41342 417832 106286
rect 418172 103514 418200 106694
rect 417896 103486 418200 103514
rect 417896 99414 417924 103486
rect 417884 99408 417936 99414
rect 417884 99350 417936 99356
rect 417792 41336 417844 41342
rect 417792 41278 417844 41284
rect 417424 35896 417476 35902
rect 417424 35838 417476 35844
rect 418816 35834 418844 129814
rect 418896 120148 418948 120154
rect 418896 120090 418948 120096
rect 418804 35828 418856 35834
rect 418804 35770 418856 35776
rect 414940 34468 414992 34474
rect 414940 34410 414992 34416
rect 418908 33046 418936 120090
rect 419000 111790 419028 186322
rect 425704 179444 425756 179450
rect 425704 179386 425756 179392
rect 424324 162920 424376 162926
rect 424324 162862 424376 162868
rect 423128 158772 423180 158778
rect 423128 158714 423180 158720
rect 423036 155984 423088 155990
rect 423036 155926 423088 155932
rect 422944 151836 422996 151842
rect 422944 151778 422996 151784
rect 421656 147688 421708 147694
rect 421656 147630 421708 147636
rect 419172 146328 419224 146334
rect 419172 146270 419224 146276
rect 419080 130280 419132 130286
rect 419080 130222 419132 130228
rect 418988 111784 419040 111790
rect 418988 111726 419040 111732
rect 418988 102196 419040 102202
rect 418988 102138 419040 102144
rect 419000 38622 419028 102138
rect 419092 57866 419120 130222
rect 419184 75886 419212 146270
rect 421564 143608 421616 143614
rect 421564 143550 421616 143556
rect 420184 130144 420236 130150
rect 420184 130086 420236 130092
rect 419172 75880 419224 75886
rect 419172 75822 419224 75828
rect 420196 60722 420224 130086
rect 420276 130076 420328 130082
rect 420276 130018 420328 130024
rect 420288 63510 420316 130018
rect 421576 74458 421604 143550
rect 421668 78674 421696 147630
rect 421932 128444 421984 128450
rect 421932 128386 421984 128392
rect 421840 111852 421892 111858
rect 421840 111794 421892 111800
rect 421748 110492 421800 110498
rect 421748 110434 421800 110440
rect 421656 78668 421708 78674
rect 421656 78610 421708 78616
rect 421564 74452 421616 74458
rect 421564 74394 421616 74400
rect 420276 63504 420328 63510
rect 420276 63446 420328 63452
rect 420184 60716 420236 60722
rect 420184 60658 420236 60664
rect 419080 57860 419132 57866
rect 419080 57802 419132 57808
rect 421760 45558 421788 110434
rect 421852 46918 421880 111794
rect 421944 92478 421972 128386
rect 421932 92472 421984 92478
rect 421932 92414 421984 92420
rect 422956 81394 422984 151778
rect 423048 85542 423076 155926
rect 423140 88262 423168 158714
rect 423220 116000 423272 116006
rect 423220 115942 423272 115948
rect 423128 88256 423180 88262
rect 423128 88198 423180 88204
rect 423036 85536 423088 85542
rect 423036 85478 423088 85484
rect 422944 81388 422996 81394
rect 422944 81330 422996 81336
rect 423232 49706 423260 115942
rect 424336 91050 424364 162862
rect 424416 161492 424468 161498
rect 424416 161434 424468 161440
rect 424324 91044 424376 91050
rect 424324 90986 424376 90992
rect 424428 89690 424456 161434
rect 424508 132524 424560 132530
rect 424508 132466 424560 132472
rect 424416 89684 424468 89690
rect 424416 89626 424468 89632
rect 424520 64870 424548 132466
rect 424600 128512 424652 128518
rect 424600 128454 424652 128460
rect 424508 64864 424560 64870
rect 424508 64806 424560 64812
rect 424612 62082 424640 128454
rect 424692 118720 424744 118726
rect 424692 118662 424744 118668
rect 424600 62076 424652 62082
rect 424600 62018 424652 62024
rect 424704 53786 424732 118662
rect 424968 108112 425020 108118
rect 424968 108054 425020 108060
rect 424980 106758 425008 108054
rect 424968 106752 425020 106758
rect 424968 106694 425020 106700
rect 425716 106282 425744 179386
rect 425796 164280 425848 164286
rect 425796 164222 425848 164228
rect 425704 106276 425756 106282
rect 425704 106218 425756 106224
rect 425808 93838 425836 164222
rect 425888 157412 425940 157418
rect 425888 157354 425940 157360
rect 425796 93832 425848 93838
rect 425796 93774 425848 93780
rect 425900 86902 425928 157354
rect 426072 138032 426124 138038
rect 426072 137974 426124 137980
rect 425980 136672 426032 136678
rect 425980 136614 426032 136620
rect 425888 86896 425940 86902
rect 425888 86838 425940 86844
rect 425992 67522 426020 136614
rect 426084 70378 426112 137974
rect 428476 114510 428504 189042
rect 428556 187740 428608 187746
rect 428556 187682 428608 187688
rect 428464 114504 428516 114510
rect 428464 114446 428516 114452
rect 428568 113150 428596 187682
rect 428648 183592 428700 183598
rect 428648 183534 428700 183540
rect 428556 113144 428608 113150
rect 428556 113086 428608 113092
rect 427820 110424 427872 110430
rect 427820 110366 427872 110372
rect 427832 108118 427860 110366
rect 428660 110362 428688 183534
rect 436744 182232 436796 182238
rect 436744 182174 436796 182180
rect 435364 178084 435416 178090
rect 435364 178026 435416 178032
rect 432604 172576 432656 172582
rect 432604 172518 432656 172524
rect 431224 171148 431276 171154
rect 431224 171090 431276 171096
rect 429844 168428 429896 168434
rect 429844 168370 429896 168376
rect 428740 167068 428792 167074
rect 428740 167010 428792 167016
rect 428648 110356 428700 110362
rect 428648 110298 428700 110304
rect 427820 108112 427872 108118
rect 427820 108054 427872 108060
rect 428752 95198 428780 167010
rect 429856 96626 429884 168370
rect 429936 142180 429988 142186
rect 429936 142122 429988 142128
rect 429844 96620 429896 96626
rect 429844 96562 429896 96568
rect 428740 95192 428792 95198
rect 428740 95134 428792 95140
rect 429948 73166 429976 142122
rect 431236 97986 431264 171090
rect 431316 135312 431368 135318
rect 431316 135254 431368 135260
rect 431224 97980 431276 97986
rect 431224 97922 431276 97928
rect 429936 73160 429988 73166
rect 429936 73102 429988 73108
rect 426072 70372 426124 70378
rect 426072 70314 426124 70320
rect 425980 67516 426032 67522
rect 425980 67458 426032 67464
rect 431328 66230 431356 135254
rect 431960 115252 432012 115258
rect 431960 115194 432012 115200
rect 431972 111874 432000 115194
rect 431880 111846 432000 111874
rect 431880 110498 431908 111846
rect 431868 110492 431920 110498
rect 431868 110434 431920 110440
rect 432616 99346 432644 172518
rect 432696 127084 432748 127090
rect 432696 127026 432748 127032
rect 432604 99340 432656 99346
rect 432604 99282 432656 99288
rect 431316 66224 431368 66230
rect 431316 66166 431368 66172
rect 432708 59362 432736 127026
rect 434076 120216 434128 120222
rect 434076 120158 434128 120164
rect 434088 115258 434116 120158
rect 434076 115252 434128 115258
rect 434076 115194 434128 115200
rect 435376 104854 435404 178026
rect 435548 130008 435600 130014
rect 435548 129950 435600 129956
rect 435456 122868 435508 122874
rect 435456 122810 435508 122816
rect 435364 104848 435416 104854
rect 435364 104790 435416 104796
rect 435364 92540 435416 92546
rect 435364 92482 435416 92488
rect 432696 59356 432748 59362
rect 432696 59298 432748 59304
rect 424692 53780 424744 53786
rect 424692 53722 424744 53728
rect 423220 49700 423272 49706
rect 423220 49642 423272 49648
rect 421840 46912 421892 46918
rect 421840 46854 421892 46860
rect 421748 45552 421800 45558
rect 421748 45494 421800 45500
rect 418988 38616 419040 38622
rect 418988 38558 419040 38564
rect 418896 33040 418948 33046
rect 418896 32982 418948 32988
rect 435376 29170 435404 92482
rect 435468 56574 435496 122810
rect 435560 74526 435588 129950
rect 436100 124500 436152 124506
rect 436100 124442 436152 124448
rect 436112 122834 436140 124442
rect 436020 122806 436140 122834
rect 436020 120222 436048 122806
rect 436008 120216 436060 120222
rect 436008 120158 436060 120164
rect 436756 107409 436784 182174
rect 521752 131504 521804 131510
rect 521752 131446 521804 131452
rect 439688 131436 439740 131442
rect 439688 131378 439740 131384
rect 472072 131436 472124 131442
rect 472072 131378 472124 131384
rect 438124 131232 438176 131238
rect 438124 131174 438176 131180
rect 437478 128752 437534 128761
rect 437478 128687 437534 128696
rect 437492 128450 437520 128687
rect 437480 128444 437532 128450
rect 437480 128386 437532 128392
rect 437478 127120 437534 127129
rect 437478 127055 437534 127064
rect 437492 127022 437520 127055
rect 437480 127016 437532 127022
rect 437480 126958 437532 126964
rect 437478 125760 437534 125769
rect 437478 125695 437534 125704
rect 437492 125662 437520 125695
rect 437480 125656 437532 125662
rect 437480 125598 437532 125604
rect 437478 124400 437534 124409
rect 437478 124335 437534 124344
rect 437492 124234 437520 124335
rect 437480 124228 437532 124234
rect 437480 124170 437532 124176
rect 437478 121952 437534 121961
rect 437478 121887 437534 121896
rect 437492 121514 437520 121887
rect 437480 121508 437532 121514
rect 437480 121450 437532 121456
rect 437478 120456 437534 120465
rect 437478 120391 437534 120400
rect 437492 120154 437520 120391
rect 437480 120148 437532 120154
rect 437480 120090 437532 120096
rect 437572 120080 437624 120086
rect 437572 120022 437624 120028
rect 437584 119649 437612 120022
rect 437570 119640 437626 119649
rect 437570 119575 437626 119584
rect 437480 118652 437532 118658
rect 437480 118594 437532 118600
rect 437492 118153 437520 118594
rect 437478 118144 437534 118153
rect 437478 118079 437534 118088
rect 436836 117360 436888 117366
rect 436836 117302 436888 117308
rect 436742 107400 436798 107409
rect 436742 107335 436798 107344
rect 435548 74520 435600 74526
rect 435548 74462 435600 74468
rect 435456 56568 435508 56574
rect 435456 56510 435508 56516
rect 436848 50833 436876 117302
rect 437480 115932 437532 115938
rect 437480 115874 437532 115880
rect 437492 115705 437520 115874
rect 437478 115696 437534 115705
rect 437478 115631 437534 115640
rect 437480 114504 437532 114510
rect 437478 114472 437480 114481
rect 437532 114472 437534 114481
rect 437478 114407 437534 114416
rect 437480 113144 437532 113150
rect 437480 113086 437532 113092
rect 437492 112849 437520 113086
rect 437478 112840 437534 112849
rect 437478 112775 437534 112784
rect 437480 111784 437532 111790
rect 437480 111726 437532 111732
rect 437492 111353 437520 111726
rect 437478 111344 437534 111353
rect 437478 111279 437534 111288
rect 437480 110356 437532 110362
rect 437480 110298 437532 110304
rect 437492 109721 437520 110298
rect 437478 109712 437534 109721
rect 437478 109647 437534 109656
rect 437480 106276 437532 106282
rect 437480 106218 437532 106224
rect 437492 106049 437520 106218
rect 437478 106040 437534 106049
rect 437478 105975 437534 105984
rect 437664 104848 437716 104854
rect 437662 104816 437664 104825
rect 437716 104816 437718 104825
rect 437662 104751 437718 104760
rect 437480 103488 437532 103494
rect 437480 103430 437532 103436
rect 437492 103057 437520 103430
rect 437478 103048 437534 103057
rect 437478 102983 437534 102992
rect 437480 102128 437532 102134
rect 437480 102070 437532 102076
rect 437492 101425 437520 102070
rect 437478 101416 437534 101425
rect 437478 101351 437534 101360
rect 437478 99376 437534 99385
rect 437478 99311 437480 99320
rect 437532 99311 437534 99320
rect 437480 99282 437532 99288
rect 437480 97980 437532 97986
rect 437480 97922 437532 97928
rect 437492 97753 437520 97922
rect 437478 97744 437534 97753
rect 437478 97679 437534 97688
rect 437480 96620 437532 96626
rect 437480 96562 437532 96568
rect 437492 96257 437520 96562
rect 437478 96248 437534 96257
rect 437478 96183 437534 96192
rect 437480 95192 437532 95198
rect 437480 95134 437532 95140
rect 437492 94761 437520 95134
rect 437478 94752 437534 94761
rect 437478 94687 437534 94696
rect 437480 93832 437532 93838
rect 437480 93774 437532 93780
rect 437492 93129 437520 93774
rect 437478 93120 437534 93129
rect 437478 93055 437534 93064
rect 437478 91080 437534 91089
rect 437478 91015 437480 91024
rect 437532 91015 437534 91024
rect 437480 90986 437532 90992
rect 437480 89684 437532 89690
rect 437480 89626 437532 89632
rect 437492 89593 437520 89626
rect 437478 89584 437534 89593
rect 437478 89519 437534 89528
rect 437480 88256 437532 88262
rect 437480 88198 437532 88204
rect 437492 87961 437520 88198
rect 437478 87952 437534 87961
rect 437478 87887 437534 87896
rect 437480 86896 437532 86902
rect 437480 86838 437532 86844
rect 437492 86465 437520 86838
rect 437478 86456 437534 86465
rect 437478 86391 437534 86400
rect 437480 85536 437532 85542
rect 437480 85478 437532 85484
rect 437492 84833 437520 85478
rect 437478 84824 437534 84833
rect 437478 84759 437534 84768
rect 437480 82816 437532 82822
rect 437478 82784 437480 82793
rect 437532 82784 437534 82793
rect 437478 82719 437534 82728
rect 437480 81388 437532 81394
rect 437480 81330 437532 81336
rect 437492 81297 437520 81330
rect 437478 81288 437534 81297
rect 437478 81223 437534 81232
rect 437480 80028 437532 80034
rect 437480 79970 437532 79976
rect 437492 79665 437520 79970
rect 437478 79656 437534 79665
rect 437478 79591 437534 79600
rect 437480 78668 437532 78674
rect 437480 78610 437532 78616
rect 437492 78169 437520 78610
rect 437478 78160 437534 78169
rect 437478 78095 437534 78104
rect 438136 77246 438164 131174
rect 439504 131164 439556 131170
rect 439504 131106 439556 131112
rect 438768 130416 438820 130422
rect 438768 130358 438820 130364
rect 438780 124506 438808 130358
rect 438768 124500 438820 124506
rect 438768 124442 438820 124448
rect 438308 90364 438360 90370
rect 438308 90306 438360 90312
rect 438216 82884 438268 82890
rect 438216 82826 438268 82832
rect 438124 77240 438176 77246
rect 438124 77182 438176 77188
rect 437480 75880 437532 75886
rect 437480 75822 437532 75828
rect 437492 75721 437520 75822
rect 437478 75712 437534 75721
rect 437478 75647 437534 75656
rect 437480 74452 437532 74458
rect 437480 74394 437532 74400
rect 437492 74361 437520 74394
rect 437478 74352 437534 74361
rect 437478 74287 437534 74296
rect 437480 73160 437532 73166
rect 437480 73102 437532 73108
rect 437492 72865 437520 73102
rect 437478 72856 437534 72865
rect 437478 72791 437534 72800
rect 437480 71732 437532 71738
rect 437480 71674 437532 71680
rect 437492 71369 437520 71674
rect 437478 71360 437534 71369
rect 437478 71295 437534 71304
rect 437480 70372 437532 70378
rect 437480 70314 437532 70320
rect 437492 69737 437520 70314
rect 437478 69728 437534 69737
rect 437478 69663 437534 69672
rect 437480 67516 437532 67522
rect 437480 67458 437532 67464
rect 437492 67425 437520 67458
rect 437478 67416 437534 67425
rect 437478 67351 437534 67360
rect 437480 66224 437532 66230
rect 437478 66192 437480 66201
rect 437532 66192 437534 66201
rect 437478 66127 437534 66136
rect 437480 64864 437532 64870
rect 437480 64806 437532 64812
rect 437492 64569 437520 64806
rect 437478 64560 437534 64569
rect 437478 64495 437534 64504
rect 437480 62076 437532 62082
rect 437480 62018 437532 62024
rect 437492 61441 437520 62018
rect 437478 61432 437534 61441
rect 437478 61367 437534 61376
rect 437480 59356 437532 59362
rect 437480 59298 437532 59304
rect 437492 59129 437520 59298
rect 437478 59120 437534 59129
rect 437478 59055 437534 59064
rect 437480 57928 437532 57934
rect 437478 57896 437480 57905
rect 437532 57896 437534 57905
rect 437478 57831 437534 57840
rect 437756 56568 437808 56574
rect 437756 56510 437808 56516
rect 437768 56409 437796 56510
rect 437754 56400 437810 56409
rect 437754 56335 437810 56344
rect 437480 55208 437532 55214
rect 437480 55150 437532 55156
rect 437492 54777 437520 55150
rect 437478 54768 437534 54777
rect 437478 54703 437534 54712
rect 437480 53780 437532 53786
rect 437480 53722 437532 53728
rect 437492 53145 437520 53722
rect 437478 53136 437534 53145
rect 437478 53071 437534 53080
rect 436834 50824 436890 50833
rect 436834 50759 436890 50768
rect 437480 49700 437532 49706
rect 437480 49642 437532 49648
rect 437492 49609 437520 49642
rect 437478 49600 437534 49609
rect 437478 49535 437534 49544
rect 437480 48272 437532 48278
rect 437480 48214 437532 48220
rect 437492 47977 437520 48214
rect 437478 47968 437534 47977
rect 437478 47903 437534 47912
rect 437480 46912 437532 46918
rect 437480 46854 437532 46860
rect 437492 46481 437520 46854
rect 437478 46472 437534 46481
rect 437478 46407 437534 46416
rect 437480 45552 437532 45558
rect 437480 45494 437532 45500
rect 437492 44849 437520 45494
rect 437478 44840 437534 44849
rect 437478 44775 437534 44784
rect 437480 42764 437532 42770
rect 437480 42706 437532 42712
rect 437492 42673 437520 42706
rect 437478 42664 437534 42673
rect 437478 42599 437534 42608
rect 437480 41336 437532 41342
rect 437478 41304 437480 41313
rect 437532 41304 437534 41313
rect 437478 41239 437534 41248
rect 437480 40044 437532 40050
rect 437480 39986 437532 39992
rect 437492 39681 437520 39986
rect 437478 39672 437534 39681
rect 437478 39607 437534 39616
rect 437480 38616 437532 38622
rect 437480 38558 437532 38564
rect 437492 38185 437520 38558
rect 437478 38176 437534 38185
rect 437478 38111 437534 38120
rect 437480 35896 437532 35902
rect 437480 35838 437532 35844
rect 437492 35737 437520 35838
rect 437478 35728 437534 35737
rect 437478 35663 437534 35672
rect 437480 34468 437532 34474
rect 437480 34410 437532 34416
rect 437492 34377 437520 34410
rect 437478 34368 437534 34377
rect 437478 34303 437534 34312
rect 437480 33108 437532 33114
rect 437480 33050 437532 33056
rect 437492 33017 437520 33050
rect 437478 33008 437534 33017
rect 437478 32943 437534 32952
rect 437480 31544 437532 31550
rect 437480 31486 437532 31492
rect 437492 31249 437520 31486
rect 437478 31240 437534 31249
rect 437478 31175 437534 31184
rect 438228 29238 438256 82826
rect 438320 63073 438348 90306
rect 438306 63064 438362 63073
rect 438306 62999 438362 63008
rect 438216 29232 438268 29238
rect 438216 29174 438268 29180
rect 435364 29164 435416 29170
rect 435364 29106 435416 29112
rect 413560 29096 413612 29102
rect 413560 29038 413612 29044
rect 439516 28898 439544 131106
rect 439596 130348 439648 130354
rect 439596 130290 439648 130296
rect 439608 37262 439636 130290
rect 439700 41410 439728 131378
rect 443184 131164 443236 131170
rect 443184 131106 443236 131112
rect 439872 130484 439924 130490
rect 439872 130426 439924 130432
rect 439780 130212 439832 130218
rect 439780 130154 439832 130160
rect 439792 67590 439820 130154
rect 439884 86970 439912 130426
rect 443196 129962 443224 131106
rect 450268 130416 450320 130422
rect 450268 130358 450320 130364
rect 450280 129962 450308 130358
rect 464528 130348 464580 130354
rect 464528 130290 464580 130296
rect 464540 129962 464568 130290
rect 439964 129940 440016 129946
rect 443196 129934 443532 129962
rect 450280 129934 450616 129962
rect 464540 129934 464876 129962
rect 439964 129882 440016 129888
rect 439976 88330 440004 129882
rect 457444 129872 457496 129878
rect 472084 129826 472112 131378
rect 478880 131368 478932 131374
rect 478880 131310 478932 131316
rect 478892 129962 478920 131310
rect 485964 131300 486016 131306
rect 485964 131242 486016 131248
rect 485976 129962 486004 131242
rect 493140 130280 493192 130286
rect 493140 130222 493192 130228
rect 493152 129962 493180 130222
rect 514898 130212 514950 130218
rect 514898 130154 514950 130160
rect 500638 130144 500690 130150
rect 500638 130086 500690 130092
rect 478892 129934 479228 129962
rect 485976 129934 486312 129962
rect 493152 129934 493488 129962
rect 500650 129948 500678 130086
rect 507400 130076 507452 130082
rect 507400 130018 507452 130024
rect 507412 129962 507440 130018
rect 507412 129934 507748 129962
rect 514910 129948 514938 130154
rect 521764 129962 521792 131446
rect 536012 131232 536064 131238
rect 536012 131174 536064 131180
rect 528836 130008 528888 130014
rect 521764 129934 522100 129962
rect 536024 129962 536052 131174
rect 528888 129956 529184 129962
rect 528836 129950 529184 129956
rect 528848 129934 529184 129950
rect 536024 129934 536360 129962
rect 539324 129940 539376 129946
rect 539324 129882 539376 129888
rect 457496 129820 457792 129826
rect 457444 129814 457792 129820
rect 457456 129798 457792 129814
rect 472052 129798 472112 129826
rect 539336 126041 539364 129882
rect 539322 126032 539378 126041
rect 539322 125967 539378 125976
rect 439964 88324 440016 88330
rect 439964 88266 440016 88272
rect 439872 86964 439924 86970
rect 439872 86906 439924 86912
rect 439872 67652 439924 67658
rect 439872 67594 439924 67600
rect 439780 67584 439832 67590
rect 439780 67526 439832 67532
rect 439780 60784 439832 60790
rect 439780 60726 439832 60732
rect 439688 41404 439740 41410
rect 439688 41346 439740 41352
rect 439596 37256 439648 37262
rect 439596 37198 439648 37204
rect 439792 30326 439820 60726
rect 439780 30320 439832 30326
rect 439780 30262 439832 30268
rect 439884 30258 439912 67594
rect 439964 55276 440016 55282
rect 439964 55218 440016 55224
rect 439872 30252 439924 30258
rect 439872 30194 439924 30200
rect 439504 28892 439556 28898
rect 439504 28834 439556 28840
rect 413468 28824 413520 28830
rect 413468 28766 413520 28772
rect 411260 28688 411312 28694
rect 411260 28630 411312 28636
rect 439976 28626 440004 55218
rect 440056 45620 440108 45626
rect 440056 45562 440108 45568
rect 440068 29306 440096 45562
rect 445004 30110 445340 30138
rect 454940 30110 455276 30138
rect 440056 29300 440108 29306
rect 440056 29242 440108 29248
rect 445312 28898 445340 30110
rect 445300 28892 445352 28898
rect 445300 28834 445352 28840
rect 455248 28762 455276 30110
rect 464632 30110 464968 30138
rect 474752 30110 474996 30138
rect 484596 30110 484932 30138
rect 494624 30110 494960 30138
rect 504652 30110 504988 30138
rect 514772 30110 514924 30138
rect 524616 30110 524952 30138
rect 534644 30110 534980 30138
rect 464632 28966 464660 30110
rect 464620 28960 464672 28966
rect 464620 28902 464672 28908
rect 455236 28756 455288 28762
rect 455236 28698 455288 28704
rect 474752 28694 474780 30110
rect 484596 29306 484624 30110
rect 484584 29300 484636 29306
rect 484584 29242 484636 29248
rect 474740 28688 474792 28694
rect 474740 28630 474792 28636
rect 494624 28626 494652 30110
rect 504652 28830 504680 30110
rect 514772 29102 514800 30110
rect 524616 29238 524644 30110
rect 524604 29232 524656 29238
rect 524604 29174 524656 29180
rect 534644 29170 534672 30110
rect 534632 29164 534684 29170
rect 534632 29106 534684 29112
rect 514760 29096 514812 29102
rect 514760 29038 514812 29044
rect 504640 28824 504692 28830
rect 504640 28766 504692 28772
rect 382280 28620 382332 28626
rect 382280 28562 382332 28568
rect 439964 28620 440016 28626
rect 439964 28562 440016 28568
rect 494612 28620 494664 28626
rect 494612 28562 494664 28568
rect 349160 28552 349212 28558
rect 349160 28494 349212 28500
rect 338120 28484 338172 28490
rect 338120 28426 338172 28432
rect 327080 28416 327132 28422
rect 327080 28358 327132 28364
rect 294052 28280 294104 28286
rect 294052 28222 294104 28228
rect 271972 28212 272024 28218
rect 271972 28154 272024 28160
rect 261116 28144 261168 28150
rect 261116 28086 261168 28092
rect 250076 28076 250128 28082
rect 250076 28018 250128 28024
rect 540256 20670 540284 202846
rect 540336 198756 540388 198762
rect 540336 198698 540388 198704
rect 540348 60722 540376 198698
rect 540428 197396 540480 197402
rect 540428 197338 540480 197344
rect 540440 100706 540468 197338
rect 542544 130484 542596 130490
rect 542544 130426 542596 130432
rect 542360 129804 542412 129810
rect 542360 129746 542412 129752
rect 541624 125656 541676 125662
rect 541624 125598 541676 125604
rect 540428 100700 540480 100706
rect 540428 100642 540480 100648
rect 540428 85604 540480 85610
rect 540428 85546 540480 85552
rect 540336 60716 540388 60722
rect 540336 60658 540388 60664
rect 540336 45620 540388 45626
rect 540336 45562 540388 45568
rect 540348 29034 540376 45562
rect 540336 29028 540388 29034
rect 540336 28970 540388 28976
rect 540440 28898 540468 85546
rect 540428 28892 540480 28898
rect 540428 28834 540480 28840
rect 541636 28762 541664 125598
rect 542372 98161 542400 129746
rect 542452 128376 542504 128382
rect 542452 128318 542504 128324
rect 542464 107273 542492 128318
rect 542556 116385 542584 130426
rect 542542 116376 542598 116385
rect 542542 116311 542598 116320
rect 542450 107264 542506 107273
rect 542450 107199 542506 107208
rect 542358 98152 542414 98161
rect 542358 98087 542414 98096
rect 542358 89040 542414 89049
rect 542358 88975 542414 88984
rect 542372 30258 542400 88975
rect 542450 80064 542506 80073
rect 542450 79999 542506 80008
rect 542464 30326 542492 79999
rect 542542 70952 542598 70961
rect 542542 70887 542598 70896
rect 542556 31686 542584 70887
rect 542634 61840 542690 61849
rect 542634 61775 542690 61784
rect 542544 31680 542596 31686
rect 542544 31622 542596 31628
rect 542648 31618 542676 61775
rect 542726 52728 542782 52737
rect 542726 52663 542782 52672
rect 542740 31754 542768 52663
rect 543016 43625 543044 218010
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 543096 178084 543148 178090
rect 543096 178026 543148 178032
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 543002 43616 543058 43625
rect 543002 43551 543058 43560
rect 543108 34649 543136 178026
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580184 125662 580212 125967
rect 580172 125656 580224 125662
rect 580172 125598 580224 125604
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580184 85610 580212 86119
rect 580172 85604 580224 85610
rect 580172 85546 580224 85552
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580184 45626 580212 46271
rect 580172 45620 580224 45626
rect 580172 45562 580224 45568
rect 543094 34640 543150 34649
rect 543094 34575 543150 34584
rect 542728 31748 542780 31754
rect 542728 31690 542780 31696
rect 542636 31612 542688 31618
rect 542636 31554 542688 31560
rect 542452 30320 542504 30326
rect 542452 30262 542504 30268
rect 542360 30252 542412 30258
rect 542360 30194 542412 30200
rect 541624 28756 541676 28762
rect 541624 28698 541676 28704
rect 540244 20664 540296 20670
rect 540244 20606 540296 20612
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 227720 6860 227772 6866
rect 227720 6802 227772 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 205640 4140 205692 4146
rect 205640 4082 205692 4088
rect 195244 4072 195296 4078
rect 195244 4014 195296 4020
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 572 3664 624 3670
rect 572 3606 624 3612
rect 1308 3664 1360 3670
rect 1308 3606 1360 3612
rect 584 480 612 3606
rect 1688 480 1716 3674
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 48226 334192 48282 334248
rect 47766 332968 47822 333024
rect 47674 330112 47730 330168
rect 47858 331064 47914 331120
rect 48134 325760 48190 325816
rect 48042 307264 48098 307320
rect 209686 334056 209742 334112
rect 208306 332832 208362 332888
rect 208214 331064 208270 331120
rect 49606 328434 49662 328490
rect 49514 327482 49570 327538
rect 49422 305586 49478 305642
rect 208122 327392 208178 327448
rect 207018 325760 207074 325816
rect 55862 299512 55918 299568
rect 67822 299512 67878 299568
rect 65798 298016 65854 298072
rect 67546 298016 67602 298072
rect 69294 298016 69350 298072
rect 70214 298016 70270 298072
rect 71686 298016 71742 298072
rect 73066 298016 73122 298072
rect 74446 298016 74502 298072
rect 75550 298016 75606 298072
rect 76838 298036 76894 298072
rect 76838 298016 76840 298036
rect 76840 298016 76892 298036
rect 76892 298016 76894 298036
rect 77114 298016 77170 298072
rect 78494 298016 78550 298072
rect 79874 298016 79930 298072
rect 81254 298016 81310 298072
rect 82634 298016 82690 298072
rect 84014 298016 84070 298072
rect 85486 298016 85542 298072
rect 86682 298016 86738 298072
rect 88154 298016 88210 298072
rect 89166 298016 89222 298072
rect 89534 298016 89590 298072
rect 91006 298016 91062 298072
rect 92294 298016 92350 298072
rect 93674 298016 93730 298072
rect 95054 298016 95110 298072
rect 96434 298016 96490 298072
rect 97078 298016 97134 298072
rect 97906 298016 97962 298072
rect 100666 298016 100722 298072
rect 101862 298016 101918 298072
rect 102966 298016 103022 298072
rect 103334 298016 103390 298072
rect 104254 298016 104310 298072
rect 104714 298016 104770 298072
rect 105542 298016 105598 298072
rect 106094 298016 106150 298072
rect 106646 298016 106702 298072
rect 107474 298016 107530 298072
rect 107750 298016 107806 298072
rect 108854 298016 108910 298072
rect 110326 298016 110382 298072
rect 111614 298016 111670 298072
rect 112994 298016 113050 298072
rect 114466 298016 114522 298072
rect 115846 298016 115902 298072
rect 117226 298016 117282 298072
rect 78586 297880 78642 297936
rect 79966 297880 80022 297936
rect 81346 297880 81402 297936
rect 82726 297880 82782 297936
rect 84106 297880 84162 297936
rect 85394 297880 85450 297936
rect 85302 297064 85358 297120
rect 86774 297880 86830 297936
rect 86866 297744 86922 297800
rect 88246 297880 88302 297936
rect 90914 297880 90970 297936
rect 92386 297880 92442 297936
rect 93582 297880 93638 297936
rect 93766 297744 93822 297800
rect 95146 297880 95202 297936
rect 96526 297880 96582 297936
rect 97814 297880 97870 297936
rect 100574 297880 100630 297936
rect 101954 297880 102010 297936
rect 102046 297744 102102 297800
rect 113086 297880 113142 297936
rect 131118 129684 131120 129704
rect 131120 129684 131172 129704
rect 131172 129684 131174 129704
rect 131118 129648 131174 129684
rect 131210 129104 131266 129160
rect 131302 128560 131358 128616
rect 131210 126812 131266 126848
rect 131210 126792 131212 126812
rect 131212 126792 131264 126812
rect 131264 126792 131266 126812
rect 131118 126112 131174 126168
rect 131118 125024 131174 125080
rect 131210 124480 131266 124536
rect 131118 123256 131174 123312
rect 131210 122748 131212 122768
rect 131212 122748 131264 122768
rect 131264 122748 131266 122768
rect 131210 122712 131266 122748
rect 131210 122032 131266 122088
rect 131118 121488 131174 121544
rect 131210 120944 131266 121000
rect 131118 119176 131174 119232
rect 131210 118652 131266 118688
rect 131210 118632 131212 118652
rect 131212 118632 131264 118652
rect 131264 118632 131266 118652
rect 131118 117952 131174 118008
rect 131210 117408 131266 117464
rect 131210 116864 131266 116920
rect 131118 116184 131174 116240
rect 131210 115640 131266 115696
rect 131210 115096 131266 115152
rect 131210 114436 131266 114472
rect 131210 114416 131212 114436
rect 131212 114416 131264 114436
rect 131264 114416 131266 114436
rect 131302 113872 131358 113928
rect 131118 113328 131174 113384
rect 131210 112784 131266 112840
rect 131118 112104 131174 112160
rect 131210 111016 131266 111072
rect 131210 110356 131266 110392
rect 131210 110336 131212 110356
rect 131212 110336 131264 110356
rect 131264 110336 131266 110356
rect 131118 109792 131174 109848
rect 131302 109248 131358 109304
rect 131210 108568 131266 108624
rect 131118 108024 131174 108080
rect 131210 107500 131266 107536
rect 131210 107480 131212 107500
rect 131212 107480 131264 107500
rect 131264 107480 131266 107500
rect 131118 106936 131174 106992
rect 131302 106256 131358 106312
rect 131118 105712 131174 105768
rect 131210 105168 131266 105224
rect 131210 104488 131266 104544
rect 131118 103944 131174 104000
rect 131210 103420 131266 103456
rect 131210 103400 131212 103420
rect 131212 103400 131264 103420
rect 131264 103400 131266 103420
rect 131670 102720 131726 102776
rect 131118 102176 131174 102232
rect 131210 101632 131266 101688
rect 131118 101088 131174 101144
rect 131210 99864 131266 99920
rect 131210 99340 131266 99376
rect 131210 99320 131212 99340
rect 131212 99320 131264 99340
rect 131264 99320 131266 99340
rect 131118 98640 131174 98696
rect 131486 98096 131542 98152
rect 131210 97552 131266 97608
rect 131118 97008 131174 97064
rect 131210 96328 131266 96384
rect 131118 95784 131174 95840
rect 131210 94560 131266 94616
rect 131118 94016 131174 94072
rect 131210 93472 131266 93528
rect 131118 92792 131174 92848
rect 131210 92284 131212 92304
rect 131212 92284 131264 92304
rect 131264 92284 131266 92304
rect 131210 92248 131266 92284
rect 131118 91704 131174 91760
rect 131302 91160 131358 91216
rect 131210 90480 131266 90536
rect 131118 89936 131174 89992
rect 131302 88712 131358 88768
rect 131210 88204 131212 88224
rect 131212 88204 131264 88224
rect 131264 88204 131266 88224
rect 131210 88168 131266 88204
rect 131118 87624 131174 87680
rect 131302 86944 131358 87000
rect 131210 86400 131266 86456
rect 131118 85856 131174 85912
rect 131118 84632 131174 84688
rect 131210 83544 131266 83600
rect 131118 82864 131174 82920
rect 131578 82320 131634 82376
rect 131210 81776 131266 81832
rect 131210 80552 131266 80608
rect 131210 80028 131266 80064
rect 131210 80008 131212 80028
rect 131212 80008 131264 80028
rect 131264 80008 131266 80028
rect 131118 79464 131174 79520
rect 131210 78784 131266 78840
rect 131210 78240 131266 78296
rect 131118 77696 131174 77752
rect 131302 77016 131358 77072
rect 131210 76472 131266 76528
rect 131118 75928 131174 75984
rect 131210 75248 131266 75304
rect 131118 74704 131174 74760
rect 131210 74160 131266 74216
rect 131118 73616 131174 73672
rect 131210 72972 131212 72992
rect 131212 72972 131264 72992
rect 131264 72972 131266 72992
rect 131210 72936 131266 72972
rect 131118 72392 131174 72448
rect 131210 71168 131266 71224
rect 131118 70624 131174 70680
rect 131210 70080 131266 70136
rect 131118 69400 131174 69456
rect 131118 68856 131174 68912
rect 131210 68312 131266 68368
rect 131302 67768 131358 67824
rect 131210 67088 131266 67144
rect 131118 66544 131174 66600
rect 131210 66000 131266 66056
rect 131118 65320 131174 65376
rect 131210 64812 131212 64832
rect 131212 64812 131264 64832
rect 131264 64812 131266 64832
rect 131210 64776 131266 64812
rect 131118 63688 131174 63744
rect 131210 61920 131266 61976
rect 131118 60696 131174 60752
rect 131670 59472 131726 59528
rect 131302 58384 131358 58440
rect 131210 57876 131212 57896
rect 131212 57876 131264 57896
rect 131264 57876 131266 57896
rect 131210 57840 131266 57876
rect 131210 57160 131266 57216
rect 131118 56616 131174 56672
rect 131210 55392 131266 55448
rect 131210 54848 131266 54904
rect 131302 53624 131358 53680
rect 131210 53080 131266 53136
rect 131118 52536 131174 52592
rect 131210 51312 131266 51368
rect 131210 50768 131266 50824
rect 131118 50224 131174 50280
rect 131302 49544 131358 49600
rect 131210 49000 131266 49056
rect 131118 48456 131174 48512
rect 131210 47232 131266 47288
rect 131210 46688 131266 46744
rect 131118 46144 131174 46200
rect 131210 45364 131212 45384
rect 131212 45364 131264 45384
rect 131264 45364 131266 45384
rect 131210 45328 131266 45364
rect 131118 44920 131174 44976
rect 131302 44376 131358 44432
rect 131210 43696 131266 43752
rect 131118 43152 131174 43208
rect 131210 42644 131212 42664
rect 131212 42644 131264 42664
rect 131264 42644 131266 42664
rect 131210 42608 131266 42644
rect 131118 41928 131174 41984
rect 131210 40840 131266 40896
rect 131118 40296 131174 40352
rect 131210 38564 131212 38584
rect 131212 38564 131264 38584
rect 131264 38564 131266 38584
rect 131210 38528 131266 38564
rect 131118 37848 131174 37904
rect 131486 37304 131542 37360
rect 131302 36760 131358 36816
rect 131210 36080 131266 36136
rect 131210 35536 131266 35592
rect 131118 34992 131174 35048
rect 131210 32680 131266 32736
rect 131118 32000 131174 32056
rect 131210 31456 131266 31512
rect 131302 30912 131358 30968
rect 131118 30368 131174 30424
rect 207018 307128 207074 307184
rect 207018 305496 207074 305552
rect 209594 329976 209650 330032
rect 209502 328480 209558 328536
rect 238574 299784 238630 299840
rect 229098 298288 229154 298344
rect 215850 298016 215906 298072
rect 224958 298016 225014 298072
rect 226338 298016 226394 298072
rect 227718 298016 227774 298072
rect 230478 298016 230534 298072
rect 231950 298016 232006 298072
rect 233238 298016 233294 298072
rect 234710 298016 234766 298072
rect 237194 298016 237250 298072
rect 229282 297744 229338 297800
rect 237378 297880 237434 297936
rect 237286 297744 237342 297800
rect 243082 299648 243138 299704
rect 238666 298016 238722 298072
rect 240138 298016 240194 298072
rect 241426 298016 241482 298072
rect 242898 298016 242954 298072
rect 238574 297064 238630 297120
rect 238758 297880 238814 297936
rect 240046 297064 240102 297120
rect 241518 297880 241574 297936
rect 242806 297744 242862 297800
rect 244094 298016 244150 298072
rect 244278 298016 244334 298072
rect 245566 298016 245622 298072
rect 246854 298016 246910 298072
rect 248234 298016 248290 298072
rect 249706 298016 249762 298072
rect 250994 298016 251050 298072
rect 252374 298016 252430 298072
rect 253754 298016 253810 298072
rect 255134 298016 255190 298072
rect 256514 298016 256570 298072
rect 257894 298016 257950 298072
rect 259182 298016 259238 298072
rect 260654 298016 260710 298072
rect 262034 298016 262090 298072
rect 263506 298016 263562 298072
rect 266174 298016 266230 298072
rect 273074 298016 273130 298072
rect 274546 298016 274602 298072
rect 275926 298016 275982 298072
rect 277306 298016 277362 298072
rect 243082 297880 243138 297936
rect 244186 297880 244242 297936
rect 246762 297880 246818 297936
rect 246946 297744 247002 297800
rect 248326 297880 248382 297936
rect 249614 297880 249670 297936
rect 251086 297880 251142 297936
rect 252282 297880 252338 297936
rect 252466 297744 252522 297800
rect 253846 297880 253902 297936
rect 255226 297880 255282 297936
rect 256606 297880 256662 297936
rect 257802 297880 257858 297936
rect 257986 297744 258042 297800
rect 259366 297880 259422 297936
rect 259274 297744 259330 297800
rect 260746 297880 260802 297936
rect 262126 297880 262182 297936
rect 263414 297880 263470 297936
rect 264794 296928 264850 296984
rect 264886 296792 264942 296848
rect 267646 297064 267702 297120
rect 267462 296928 267518 296984
rect 266266 296792 266322 296848
rect 267554 296792 267610 296848
rect 269026 296792 269082 296848
rect 270406 296792 270462 296848
rect 271786 296792 271842 296848
rect 273166 296792 273222 296848
rect 408958 251776 409014 251832
rect 408866 249600 408922 249656
rect 186318 249464 186374 249520
rect 186318 248276 186320 248296
rect 186320 248276 186372 248296
rect 186372 248276 186374 248296
rect 186318 248240 186374 248276
rect 186410 247152 186466 247208
rect 186318 245928 186374 245984
rect 186318 244840 186374 244896
rect 186318 243616 186374 243672
rect 186318 242528 186374 242584
rect 186318 241304 186374 241360
rect 186318 240080 186374 240136
rect 186410 238992 186466 239048
rect 409418 248240 409474 248296
rect 409326 247696 409382 247752
rect 409326 245520 409382 245576
rect 409326 243616 409382 243672
rect 409326 241576 409382 241632
rect 187146 237768 187202 237824
rect 186318 236680 186374 236736
rect 186318 235456 186374 235512
rect 186318 234368 186374 234424
rect 186318 233164 186374 233200
rect 186318 233144 186320 233164
rect 186320 233144 186372 233164
rect 186372 233144 186374 233164
rect 186410 232056 186466 232112
rect 186318 230832 186374 230888
rect 186318 229608 186374 229664
rect 186318 228520 186374 228576
rect 132222 127880 132278 127936
rect 132038 127336 132094 127392
rect 132038 125568 132094 125624
rect 132222 123800 132278 123856
rect 131946 120264 132002 120320
rect 132222 119720 132278 119776
rect 132130 111560 132186 111616
rect 131854 100408 131910 100464
rect 132222 95240 132278 95296
rect 131854 64232 131910 64288
rect 132222 89392 132278 89448
rect 131946 62464 132002 62520
rect 132222 85312 132278 85368
rect 132222 84088 132278 84144
rect 132222 81096 132278 81152
rect 132222 63008 132278 63064
rect 132130 61240 132186 61296
rect 132222 60152 132278 60208
rect 132038 58928 132094 58984
rect 132222 56072 132278 56128
rect 132498 71848 132554 71904
rect 132498 54304 132554 54360
rect 132314 51992 132370 52048
rect 131946 47776 132002 47832
rect 131854 41384 131910 41440
rect 131946 39616 132002 39672
rect 132498 39072 132554 39128
rect 131854 34448 131910 34504
rect 132130 33768 132186 33824
rect 132222 33224 132278 33280
rect 186318 227296 186374 227352
rect 186410 226208 186466 226264
rect 186318 225004 186374 225040
rect 186318 224984 186320 225004
rect 186320 224984 186372 225004
rect 186372 224984 186374 225004
rect 186318 223896 186374 223952
rect 186318 222672 186374 222728
rect 186318 221448 186374 221504
rect 186318 220360 186374 220416
rect 186410 219136 186466 219192
rect 186318 218068 186374 218104
rect 186318 218048 186320 218068
rect 186320 218048 186372 218068
rect 186372 218048 186374 218068
rect 186318 216824 186374 216880
rect 186318 215736 186374 215792
rect 186318 214512 186374 214568
rect 186318 213424 186374 213480
rect 186318 212200 186374 212256
rect 186410 210976 186466 211032
rect 186318 209908 186374 209944
rect 186318 209888 186320 209908
rect 186320 209888 186372 209908
rect 186372 209888 186374 209908
rect 186962 208664 187018 208720
rect 186318 207576 186374 207632
rect 186318 206352 186374 206408
rect 186318 205264 186374 205320
rect 186410 204040 186466 204096
rect 186318 202972 186374 203008
rect 186318 202952 186320 202972
rect 186320 202952 186372 202972
rect 186372 202952 186374 202972
rect 186318 201728 186374 201784
rect 186318 200504 186374 200560
rect 186318 199416 186374 199472
rect 186318 198192 186374 198248
rect 186410 195880 186466 195936
rect 186318 194792 186374 194848
rect 186318 193568 186374 193624
rect 186318 192344 186374 192400
rect 186318 191256 186374 191312
rect 186318 190032 186374 190088
rect 186410 188944 186466 189000
rect 186318 187740 186374 187776
rect 186318 187720 186320 187740
rect 186320 187720 186372 187740
rect 186372 187720 186374 187740
rect 186318 186632 186374 186688
rect 186318 185408 186374 185464
rect 186318 184320 186374 184376
rect 186318 183096 186374 183152
rect 186410 181872 186466 181928
rect 186318 180784 186374 180840
rect 186318 179560 186374 179616
rect 186318 178472 186374 178528
rect 186318 177248 186374 177304
rect 186318 176160 186374 176216
rect 186318 174936 186374 174992
rect 186410 173712 186466 173768
rect 186318 172644 186374 172680
rect 186318 172624 186320 172644
rect 186320 172624 186372 172644
rect 186372 172624 186374 172644
rect 186318 171400 186374 171456
rect 186318 170312 186374 170368
rect 186318 169088 186374 169144
rect 186318 168000 186374 168056
rect 186410 166776 186466 166832
rect 186318 165708 186374 165744
rect 186318 165688 186320 165708
rect 186320 165688 186372 165708
rect 186372 165688 186374 165708
rect 186318 164464 186374 164520
rect 186318 163240 186374 163296
rect 186318 162152 186374 162208
rect 186318 160928 186374 160984
rect 186318 159840 186374 159896
rect 186410 158616 186466 158672
rect 186318 157528 186374 157584
rect 186318 156304 186374 156360
rect 186318 155216 186374 155272
rect 186318 153992 186374 154048
rect 186318 152768 186374 152824
rect 186410 151680 186466 151736
rect 186318 150476 186374 150512
rect 186318 150456 186320 150476
rect 186320 150456 186372 150476
rect 186372 150456 186374 150476
rect 186318 149368 186374 149424
rect 186318 148144 186374 148200
rect 186318 147056 186374 147112
rect 186318 145832 186374 145888
rect 186410 144608 186466 144664
rect 186318 143520 186374 143576
rect 186318 142296 186374 142352
rect 186318 139984 186374 140040
rect 186318 138896 186374 138952
rect 186318 137672 186374 137728
rect 186410 136584 186466 136640
rect 186318 135360 186374 135416
rect 186318 133048 186374 133104
rect 186318 131824 186374 131880
rect 186318 130736 186374 130792
rect 186410 129512 186466 129568
rect 186318 128424 186374 128480
rect 186318 127200 186374 127256
rect 186318 125976 186374 126032
rect 186318 124888 186374 124944
rect 186318 122576 186374 122632
rect 186410 121352 186466 121408
rect 186318 120264 186374 120320
rect 409970 217232 410026 217288
rect 410246 228112 410302 228168
rect 410522 239536 410578 239592
rect 410430 231920 410486 231976
rect 410338 226208 410394 226264
rect 410154 224304 410210 224360
rect 410062 213560 410118 213616
rect 409878 209480 409934 209536
rect 411350 214784 411406 214840
rect 411626 230016 411682 230072
rect 411534 220496 411590 220552
rect 411902 235728 411958 235784
rect 411810 222400 411866 222456
rect 580170 219000 580226 219056
rect 411718 218592 411774 218648
rect 411442 211112 411498 211168
rect 411258 207304 411314 207360
rect 409326 205536 409382 205592
rect 411258 203496 411314 203552
rect 411258 201612 411314 201648
rect 411258 201592 411260 201612
rect 411260 201592 411312 201612
rect 411312 201592 411314 201612
rect 411258 199688 411314 199744
rect 411258 197784 411314 197840
rect 187054 197104 187110 197160
rect 186318 119040 186374 119096
rect 186318 117952 186374 118008
rect 186318 116728 186374 116784
rect 186318 115504 186374 115560
rect 411994 195880 412050 195936
rect 411258 193976 411314 194032
rect 411902 192072 411958 192128
rect 187146 141208 187202 141264
rect 186962 113192 187018 113248
rect 186318 112104 186374 112160
rect 186318 110880 186374 110936
rect 186318 109792 186374 109848
rect 186318 108568 186374 108624
rect 186410 107480 186466 107536
rect 186318 106292 186320 106312
rect 186320 106292 186372 106312
rect 186372 106292 186374 106312
rect 186318 106256 186374 106292
rect 186318 105032 186374 105088
rect 186318 103944 186374 104000
rect 186318 102720 186374 102776
rect 186318 101632 186374 101688
rect 186318 100408 186374 100464
rect 186410 99320 186466 99376
rect 186318 98096 186374 98152
rect 186318 96872 186374 96928
rect 186318 95784 186374 95840
rect 186318 94560 186374 94616
rect 186318 93472 186374 93528
rect 186318 91160 186374 91216
rect 186318 89936 186374 89992
rect 186318 88848 186374 88904
rect 186318 87624 186374 87680
rect 186318 86400 186374 86456
rect 186410 84088 186466 84144
rect 186318 83000 186374 83056
rect 186318 80688 186374 80744
rect 186318 79464 186374 79520
rect 186410 77152 186466 77208
rect 186318 75964 186320 75984
rect 186320 75964 186372 75984
rect 186372 75964 186374 75984
rect 186318 75928 186374 75964
rect 187238 134136 187294 134192
rect 187054 85312 187110 85368
rect 186318 73616 186374 73672
rect 186318 72528 186374 72584
rect 186318 71304 186374 71360
rect 186410 70216 186466 70272
rect 186318 69028 186320 69048
rect 186320 69028 186372 69048
rect 186372 69028 186374 69048
rect 186318 68992 186374 69028
rect 186318 67768 186374 67824
rect 186318 66680 186374 66736
rect 186318 65456 186374 65512
rect 186318 64368 186374 64424
rect 186318 63144 186374 63200
rect 186410 62056 186466 62112
rect 186318 60852 186374 60888
rect 186318 60832 186320 60852
rect 186320 60832 186372 60852
rect 186372 60832 186374 60852
rect 186318 59744 186374 59800
rect 186318 58520 186374 58576
rect 187330 123664 187386 123720
rect 187146 81776 187202 81832
rect 186962 57296 187018 57352
rect 186318 56208 186374 56264
rect 186318 54984 186374 55040
rect 186318 52672 186374 52728
rect 186318 51584 186374 51640
rect 186318 49136 186374 49192
rect 186318 48048 186374 48104
rect 186318 44512 186374 44568
rect 187422 114416 187478 114472
rect 187514 92248 187570 92304
rect 187422 78240 187478 78296
rect 187238 74840 187294 74896
rect 187054 53896 187110 53952
rect 186318 43424 186374 43480
rect 187146 50360 187202 50416
rect 186410 42200 186466 42256
rect 186318 38684 186374 38720
rect 186318 38664 186320 38684
rect 186320 38664 186372 38684
rect 186372 38664 186374 38684
rect 186318 37576 186374 37632
rect 187422 46824 187478 46880
rect 187238 45736 187294 45792
rect 186962 41112 187018 41168
rect 186318 36352 186374 36408
rect 187054 39888 187110 39944
rect 186410 35264 186466 35320
rect 186318 34040 186374 34096
rect 186410 32952 186466 33008
rect 186318 31764 186320 31784
rect 186320 31764 186372 31784
rect 186372 31764 186374 31784
rect 186318 31728 186374 31764
rect 186318 30640 186374 30696
rect 411258 190168 411314 190224
rect 411258 188264 411314 188320
rect 411258 186380 411314 186416
rect 411258 186360 411260 186380
rect 411260 186360 411312 186380
rect 411312 186360 411314 186380
rect 411258 184456 411314 184512
rect 411258 182552 411314 182608
rect 411258 180648 411314 180704
rect 411258 178744 411314 178800
rect 411258 176976 411314 177032
rect 411258 175072 411314 175128
rect 411258 173168 411314 173224
rect 411258 171264 411314 171320
rect 411258 169360 411314 169416
rect 411258 167456 411314 167512
rect 411258 165552 411314 165608
rect 411258 163648 411314 163704
rect 411258 161744 411314 161800
rect 411258 159840 411314 159896
rect 411258 157936 411314 157992
rect 411258 156032 411314 156088
rect 411258 154128 411314 154184
rect 411258 152224 411314 152280
rect 411258 150320 411314 150376
rect 411258 148416 411314 148472
rect 411258 146512 411314 146568
rect 411258 144608 411314 144664
rect 411258 142704 411314 142760
rect 411258 140936 411314 140992
rect 411258 139032 411314 139088
rect 411258 137128 411314 137184
rect 411258 135260 411260 135280
rect 411260 135260 411312 135280
rect 411312 135260 411314 135280
rect 411258 135224 411314 135260
rect 411258 133320 411314 133376
rect 411258 131416 411314 131472
rect 411258 129512 411314 129568
rect 411258 127608 411314 127664
rect 411258 125724 411314 125760
rect 411258 125704 411260 125724
rect 411260 125704 411312 125724
rect 411312 125704 411314 125724
rect 411258 123800 411314 123856
rect 411258 121896 411314 121952
rect 411258 119992 411314 120048
rect 411258 118088 411314 118144
rect 411258 116184 411314 116240
rect 411994 114280 412050 114336
rect 411258 112376 411314 112432
rect 411258 110492 411314 110528
rect 411258 110472 411260 110492
rect 411260 110472 411312 110492
rect 411312 110472 411314 110492
rect 411902 108568 411958 108624
rect 411258 106664 411314 106720
rect 411258 104760 411314 104816
rect 411258 102992 411314 103048
rect 411258 101088 411314 101144
rect 411258 99184 411314 99240
rect 411810 95376 411866 95432
rect 411350 93472 411406 93528
rect 411258 91568 411314 91624
rect 411258 89684 411314 89720
rect 411258 89664 411260 89684
rect 411260 89664 411312 89684
rect 411312 89664 411314 89684
rect 411258 87760 411314 87816
rect 411258 85856 411314 85912
rect 411258 83952 411314 84008
rect 411258 80164 411314 80200
rect 411258 80144 411260 80164
rect 411260 80144 411312 80164
rect 411312 80144 411314 80164
rect 411258 78276 411260 78296
rect 411260 78276 411312 78296
rect 411312 78276 411314 78296
rect 411258 78240 411314 78276
rect 411258 76336 411314 76392
rect 411258 74468 411260 74488
rect 411260 74468 411312 74488
rect 411312 74468 411314 74488
rect 411258 74432 411314 74468
rect 411258 72528 411314 72584
rect 411350 68720 411406 68776
rect 411258 66952 411314 67008
rect 411258 65068 411314 65104
rect 411258 65048 411260 65068
rect 411260 65048 411312 65068
rect 411312 65048 411314 65068
rect 411258 63144 411314 63200
rect 411258 61240 411314 61296
rect 411350 59336 411406 59392
rect 411258 57432 411314 57488
rect 411258 55528 411314 55584
rect 411258 49816 411314 49872
rect 411258 47912 411314 47968
rect 411258 46008 411314 46064
rect 411810 44104 411866 44160
rect 411258 42200 411314 42256
rect 411258 40296 411314 40352
rect 411258 38392 411314 38448
rect 411258 36488 411314 36544
rect 411258 34584 411314 34640
rect 411258 32680 411314 32736
rect 412086 97280 412142 97336
rect 412454 82048 412510 82104
rect 412362 70624 412418 70680
rect 412270 53624 412326 53680
rect 412362 51720 412418 51776
rect 411258 30912 411314 30968
rect 437478 128696 437534 128752
rect 437478 127064 437534 127120
rect 437478 125704 437534 125760
rect 437478 124344 437534 124400
rect 437478 121896 437534 121952
rect 437478 120400 437534 120456
rect 437570 119584 437626 119640
rect 437478 118088 437534 118144
rect 436742 107344 436798 107400
rect 437478 115640 437534 115696
rect 437478 114452 437480 114472
rect 437480 114452 437532 114472
rect 437532 114452 437534 114472
rect 437478 114416 437534 114452
rect 437478 112784 437534 112840
rect 437478 111288 437534 111344
rect 437478 109656 437534 109712
rect 437478 105984 437534 106040
rect 437662 104796 437664 104816
rect 437664 104796 437716 104816
rect 437716 104796 437718 104816
rect 437662 104760 437718 104796
rect 437478 102992 437534 103048
rect 437478 101360 437534 101416
rect 437478 99340 437534 99376
rect 437478 99320 437480 99340
rect 437480 99320 437532 99340
rect 437532 99320 437534 99340
rect 437478 97688 437534 97744
rect 437478 96192 437534 96248
rect 437478 94696 437534 94752
rect 437478 93064 437534 93120
rect 437478 91044 437534 91080
rect 437478 91024 437480 91044
rect 437480 91024 437532 91044
rect 437532 91024 437534 91044
rect 437478 89528 437534 89584
rect 437478 87896 437534 87952
rect 437478 86400 437534 86456
rect 437478 84768 437534 84824
rect 437478 82764 437480 82784
rect 437480 82764 437532 82784
rect 437532 82764 437534 82784
rect 437478 82728 437534 82764
rect 437478 81232 437534 81288
rect 437478 79600 437534 79656
rect 437478 78104 437534 78160
rect 437478 75656 437534 75712
rect 437478 74296 437534 74352
rect 437478 72800 437534 72856
rect 437478 71304 437534 71360
rect 437478 69672 437534 69728
rect 437478 67360 437534 67416
rect 437478 66172 437480 66192
rect 437480 66172 437532 66192
rect 437532 66172 437534 66192
rect 437478 66136 437534 66172
rect 437478 64504 437534 64560
rect 437478 61376 437534 61432
rect 437478 59064 437534 59120
rect 437478 57876 437480 57896
rect 437480 57876 437532 57896
rect 437532 57876 437534 57896
rect 437478 57840 437534 57876
rect 437754 56344 437810 56400
rect 437478 54712 437534 54768
rect 437478 53080 437534 53136
rect 436834 50768 436890 50824
rect 437478 49544 437534 49600
rect 437478 47912 437534 47968
rect 437478 46416 437534 46472
rect 437478 44784 437534 44840
rect 437478 42608 437534 42664
rect 437478 41284 437480 41304
rect 437480 41284 437532 41304
rect 437532 41284 437534 41304
rect 437478 41248 437534 41284
rect 437478 39616 437534 39672
rect 437478 38120 437534 38176
rect 437478 35672 437534 35728
rect 437478 34312 437534 34368
rect 437478 32952 437534 33008
rect 437478 31184 437534 31240
rect 438306 63008 438362 63064
rect 539322 125976 539378 126032
rect 542542 116320 542598 116376
rect 542450 107208 542506 107264
rect 542358 98096 542414 98152
rect 542358 88984 542414 89040
rect 542450 80008 542506 80064
rect 542542 70896 542598 70952
rect 542634 61784 542690 61840
rect 542726 52672 542782 52728
rect 580170 179152 580226 179208
rect 543002 43560 543058 43616
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 543094 34584 543150 34640
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect 48221 334250 48287 334253
rect 48221 334248 49434 334250
rect 48221 334192 48226 334248
rect 48282 334204 49434 334248
rect 48282 334192 50048 334204
rect 48221 334190 50048 334192
rect 48221 334187 48287 334190
rect 49374 334144 50048 334190
rect 209730 334144 210032 334204
rect 209730 334117 209790 334144
rect 209681 334112 209790 334117
rect 209681 334056 209686 334112
rect 209742 334056 209790 334112
rect 209681 334054 209790 334056
rect 209681 334051 209747 334054
rect 47761 333026 47827 333029
rect 47761 333024 49434 333026
rect 47761 332968 47766 333024
rect 47822 332980 49434 333024
rect 47822 332968 50048 332980
rect 47761 332966 50048 332968
rect 47761 332963 47827 332966
rect 49374 332920 50048 332966
rect 209730 332920 210032 332980
rect 208301 332890 208367 332893
rect 209730 332890 209790 332920
rect 208301 332888 209790 332890
rect 208301 332832 208306 332888
rect 208362 332832 209790 332888
rect 208301 332830 209790 332832
rect 208301 332827 208367 332830
rect -960 332196 480 332436
rect 49742 331152 50048 331212
rect 209730 331152 210032 331212
rect 47853 331122 47919 331125
rect 49742 331122 49802 331152
rect 47853 331120 49802 331122
rect 47853 331064 47858 331120
rect 47914 331064 49802 331120
rect 47853 331062 49802 331064
rect 208209 331122 208275 331125
rect 209730 331122 209790 331152
rect 208209 331120 209790 331122
rect 208209 331064 208214 331120
rect 208270 331064 209790 331120
rect 208209 331062 209790 331064
rect 47853 331059 47919 331062
rect 208209 331059 208275 331062
rect 47669 330170 47735 330173
rect 47669 330168 49434 330170
rect 47669 330112 47674 330168
rect 47730 330124 49434 330168
rect 47730 330112 50048 330124
rect 47669 330110 50048 330112
rect 47669 330107 47735 330110
rect 49374 330064 50048 330110
rect 209730 330064 210032 330124
rect 209589 330034 209655 330037
rect 209730 330034 209790 330064
rect 209589 330032 209790 330034
rect 209589 329976 209594 330032
rect 209650 329976 209790 330032
rect 209589 329974 209790 329976
rect 209589 329971 209655 329974
rect 209497 328538 209563 328541
rect 209497 328536 209790 328538
rect 49601 328492 49667 328495
rect 49601 328490 50048 328492
rect 49601 328434 49606 328490
rect 49662 328434 50048 328490
rect 209497 328480 209502 328536
rect 209558 328492 209790 328536
rect 209558 328480 210032 328492
rect 209497 328478 210032 328480
rect 209497 328475 209563 328478
rect 49601 328432 50048 328434
rect 209730 328432 210032 328478
rect 49601 328429 49667 328432
rect 49509 327540 49575 327543
rect 49509 327538 50048 327540
rect 49509 327482 49514 327538
rect 49570 327482 50048 327538
rect 49509 327480 50048 327482
rect 209730 327480 210032 327540
rect 49509 327477 49575 327480
rect 208117 327450 208183 327453
rect 209730 327450 209790 327480
rect 208117 327448 209790 327450
rect 208117 327392 208122 327448
rect 208178 327392 209790 327448
rect 208117 327390 209790 327392
rect 208117 327387 208183 327390
rect 48129 325818 48195 325821
rect 207013 325818 207079 325821
rect 48129 325816 49434 325818
rect 48129 325760 48134 325816
rect 48190 325772 49434 325816
rect 207013 325816 209790 325818
rect 48190 325760 50048 325772
rect 48129 325758 50048 325760
rect 48129 325755 48195 325758
rect 49374 325712 50048 325758
rect 207013 325760 207018 325816
rect 207074 325772 209790 325816
rect 207074 325760 210032 325772
rect 207013 325758 210032 325760
rect 207013 325755 207079 325758
rect 209730 325712 210032 325758
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect 48037 307322 48103 307325
rect 48037 307320 49434 307322
rect 48037 307264 48042 307320
rect 48098 307276 49434 307320
rect 48098 307264 50048 307276
rect 48037 307262 50048 307264
rect 48037 307259 48103 307262
rect 49374 307216 50048 307262
rect 209730 307216 210032 307276
rect 207013 307186 207079 307189
rect 209730 307186 209790 307216
rect 207013 307184 209790 307186
rect 207013 307128 207018 307184
rect 207074 307128 209790 307184
rect 207013 307126 209790 307128
rect 207013 307123 207079 307126
rect -960 306084 480 306324
rect 49417 305644 49483 305647
rect 49417 305642 50048 305644
rect 49417 305586 49422 305642
rect 49478 305586 50048 305642
rect 49417 305584 50048 305586
rect 209730 305584 210032 305644
rect 49417 305581 49483 305584
rect 207013 305554 207079 305557
rect 209730 305554 209790 305584
rect 207013 305552 209790 305554
rect 207013 305496 207018 305552
rect 207074 305496 209790 305552
rect 207013 305494 209790 305496
rect 207013 305491 207079 305494
rect 238569 299842 238635 299845
rect 239648 299842 239654 299844
rect 238569 299840 239654 299842
rect 238569 299784 238574 299840
rect 238630 299784 239654 299840
rect 238569 299782 239654 299784
rect 238569 299779 238635 299782
rect 239648 299780 239654 299782
rect 239718 299780 239724 299844
rect 243077 299708 243143 299709
rect 243048 299706 243054 299708
rect 242986 299646 243054 299706
rect 243118 299704 243143 299708
rect 243138 299648 243143 299704
rect 243048 299644 243054 299646
rect 243118 299644 243143 299648
rect 243077 299643 243143 299644
rect 55857 299572 55923 299573
rect 67817 299572 67883 299573
rect 55848 299570 55854 299572
rect 55766 299510 55854 299570
rect 55848 299508 55854 299510
rect 55918 299508 55924 299572
rect 67816 299508 67822 299572
rect 67886 299570 67892 299572
rect 67886 299510 67974 299570
rect 67886 299508 67892 299510
rect 55857 299507 55923 299508
rect 67817 299507 67883 299508
rect 583520 298604 584960 298844
rect 229093 298348 229159 298349
rect 229093 298344 229140 298348
rect 229204 298346 229210 298348
rect 229093 298288 229098 298344
rect 229093 298284 229140 298288
rect 229204 298286 229250 298346
rect 229204 298284 229210 298286
rect 229093 298283 229159 298284
rect 73654 298148 73660 298212
rect 73724 298148 73730 298212
rect 77886 298148 77892 298212
rect 77956 298148 77962 298212
rect 81750 298148 81756 298212
rect 81820 298148 81826 298212
rect 85430 298148 85436 298212
rect 85500 298148 85506 298212
rect 91870 298148 91876 298212
rect 91940 298148 91946 298212
rect 95550 298148 95556 298212
rect 95620 298148 95626 298212
rect 95918 298148 95924 298212
rect 95988 298148 95994 298212
rect 99414 298148 99420 298212
rect 99484 298148 99490 298212
rect 102910 298148 102916 298212
rect 102980 298148 102986 298212
rect 103278 298148 103284 298212
rect 103348 298148 103354 298212
rect 225454 298148 225460 298212
rect 225524 298148 225530 298212
rect 257838 298148 257844 298212
rect 257908 298148 257914 298212
rect 261518 298148 261524 298212
rect 261588 298148 261594 298212
rect 261886 298148 261892 298212
rect 261956 298148 261962 298212
rect 265198 298148 265204 298212
rect 265268 298148 265274 298212
rect 271822 298148 271828 298212
rect 271892 298148 271898 298212
rect 275502 298148 275508 298212
rect 275572 298148 275578 298212
rect 65558 298012 65564 298076
rect 65628 298074 65634 298076
rect 65793 298074 65859 298077
rect 65628 298072 65859 298074
rect 65628 298016 65798 298072
rect 65854 298016 65859 298072
rect 65628 298014 65859 298016
rect 65628 298012 65634 298014
rect 65793 298011 65859 298014
rect 66662 298012 66668 298076
rect 66732 298074 66738 298076
rect 67541 298074 67607 298077
rect 69289 298076 69355 298077
rect 70209 298076 70275 298077
rect 69238 298074 69244 298076
rect 66732 298072 67607 298074
rect 66732 298016 67546 298072
rect 67602 298016 67607 298072
rect 66732 298014 67607 298016
rect 69198 298014 69244 298074
rect 69308 298072 69355 298076
rect 70158 298074 70164 298076
rect 69350 298016 69355 298072
rect 66732 298012 66738 298014
rect 67541 298011 67607 298014
rect 69238 298012 69244 298014
rect 69308 298012 69355 298016
rect 70118 298014 70164 298074
rect 70228 298072 70275 298076
rect 70270 298016 70275 298072
rect 70158 298012 70164 298014
rect 70228 298012 70275 298016
rect 71446 298012 71452 298076
rect 71516 298074 71522 298076
rect 71681 298074 71747 298077
rect 71516 298072 71747 298074
rect 71516 298016 71686 298072
rect 71742 298016 71747 298072
rect 71516 298014 71747 298016
rect 71516 298012 71522 298014
rect 69289 298011 69355 298012
rect 70209 298011 70275 298012
rect 71681 298011 71747 298014
rect 72550 298012 72556 298076
rect 72620 298074 72626 298076
rect 73061 298074 73127 298077
rect 72620 298072 73127 298074
rect 72620 298016 73066 298072
rect 73122 298016 73127 298072
rect 72620 298014 73127 298016
rect 73662 298074 73722 298148
rect 74441 298074 74507 298077
rect 73662 298072 74507 298074
rect 73662 298016 74446 298072
rect 74502 298016 74507 298072
rect 73662 298014 74507 298016
rect 72620 298012 72626 298014
rect 73061 298011 73127 298014
rect 74441 298011 74507 298014
rect 75126 298012 75132 298076
rect 75196 298074 75202 298076
rect 75545 298074 75611 298077
rect 75196 298072 75611 298074
rect 75196 298016 75550 298072
rect 75606 298016 75611 298072
rect 75196 298014 75611 298016
rect 75196 298012 75202 298014
rect 75545 298011 75611 298014
rect 76230 298012 76236 298076
rect 76300 298074 76306 298076
rect 76833 298074 76899 298077
rect 76300 298072 76899 298074
rect 76300 298016 76838 298072
rect 76894 298016 76899 298072
rect 76300 298014 76899 298016
rect 76300 298012 76306 298014
rect 76833 298011 76899 298014
rect 77109 298076 77175 298077
rect 77109 298072 77156 298076
rect 77220 298074 77226 298076
rect 77109 298016 77114 298072
rect 77109 298012 77156 298016
rect 77220 298014 77266 298074
rect 77220 298012 77226 298014
rect 77109 298011 77175 298012
rect 77894 297938 77954 298148
rect 78254 298012 78260 298076
rect 78324 298074 78330 298076
rect 78489 298074 78555 298077
rect 78324 298072 78555 298074
rect 78324 298016 78494 298072
rect 78550 298016 78555 298072
rect 78324 298014 78555 298016
rect 78324 298012 78330 298014
rect 78489 298011 78555 298014
rect 79726 298012 79732 298076
rect 79796 298074 79802 298076
rect 79869 298074 79935 298077
rect 79796 298072 79935 298074
rect 79796 298016 79874 298072
rect 79930 298016 79935 298072
rect 79796 298014 79935 298016
rect 79796 298012 79802 298014
rect 79869 298011 79935 298014
rect 80830 298012 80836 298076
rect 80900 298074 80906 298076
rect 81249 298074 81315 298077
rect 80900 298072 81315 298074
rect 80900 298016 81254 298072
rect 81310 298016 81315 298072
rect 80900 298014 81315 298016
rect 80900 298012 80906 298014
rect 81249 298011 81315 298014
rect 78581 297938 78647 297941
rect 77894 297936 78647 297938
rect 77894 297880 78586 297936
rect 78642 297880 78647 297936
rect 77894 297878 78647 297880
rect 78581 297875 78647 297878
rect 79358 297876 79364 297940
rect 79428 297938 79434 297940
rect 79961 297938 80027 297941
rect 79428 297936 80027 297938
rect 79428 297880 79966 297936
rect 80022 297880 80027 297936
rect 79428 297878 80027 297880
rect 79428 297876 79434 297878
rect 79961 297875 80027 297878
rect 80278 297876 80284 297940
rect 80348 297938 80354 297940
rect 81341 297938 81407 297941
rect 80348 297936 81407 297938
rect 80348 297880 81346 297936
rect 81402 297880 81407 297936
rect 80348 297878 81407 297880
rect 81758 297938 81818 298148
rect 85438 298077 85498 298148
rect 82118 298012 82124 298076
rect 82188 298074 82194 298076
rect 82629 298074 82695 298077
rect 82188 298072 82695 298074
rect 82188 298016 82634 298072
rect 82690 298016 82695 298072
rect 82188 298014 82695 298016
rect 82188 298012 82194 298014
rect 82629 298011 82695 298014
rect 83222 298012 83228 298076
rect 83292 298074 83298 298076
rect 84009 298074 84075 298077
rect 83292 298072 84075 298074
rect 83292 298016 84014 298072
rect 84070 298016 84075 298072
rect 83292 298014 84075 298016
rect 85438 298072 85547 298077
rect 85438 298016 85486 298072
rect 85542 298016 85547 298072
rect 85438 298014 85547 298016
rect 83292 298012 83298 298014
rect 84009 298011 84075 298014
rect 85481 298011 85547 298014
rect 86534 298012 86540 298076
rect 86604 298074 86610 298076
rect 86677 298074 86743 298077
rect 86604 298072 86743 298074
rect 86604 298016 86682 298072
rect 86738 298016 86743 298072
rect 86604 298014 86743 298016
rect 86604 298012 86610 298014
rect 86677 298011 86743 298014
rect 87822 298012 87828 298076
rect 87892 298074 87898 298076
rect 88149 298074 88215 298077
rect 87892 298072 88215 298074
rect 87892 298016 88154 298072
rect 88210 298016 88215 298072
rect 87892 298014 88215 298016
rect 87892 298012 87898 298014
rect 88149 298011 88215 298014
rect 88926 298012 88932 298076
rect 88996 298074 89002 298076
rect 89161 298074 89227 298077
rect 88996 298072 89227 298074
rect 88996 298016 89166 298072
rect 89222 298016 89227 298072
rect 88996 298014 89227 298016
rect 88996 298012 89002 298014
rect 89161 298011 89227 298014
rect 89294 298012 89300 298076
rect 89364 298074 89370 298076
rect 89529 298074 89595 298077
rect 89364 298072 89595 298074
rect 89364 298016 89534 298072
rect 89590 298016 89595 298072
rect 89364 298014 89595 298016
rect 89364 298012 89370 298014
rect 89529 298011 89595 298014
rect 90766 298012 90772 298076
rect 90836 298074 90842 298076
rect 91001 298074 91067 298077
rect 90836 298072 91067 298074
rect 90836 298016 91006 298072
rect 91062 298016 91067 298072
rect 90836 298014 91067 298016
rect 91878 298074 91938 298148
rect 92289 298074 92355 298077
rect 91878 298072 92355 298074
rect 91878 298016 92294 298072
rect 92350 298016 92355 298072
rect 91878 298014 92355 298016
rect 90836 298012 90842 298014
rect 91001 298011 91067 298014
rect 92289 298011 92355 298014
rect 93526 298012 93532 298076
rect 93596 298074 93602 298076
rect 93669 298074 93735 298077
rect 95049 298076 95115 298077
rect 94998 298074 95004 298076
rect 93596 298072 93735 298074
rect 93596 298016 93674 298072
rect 93730 298016 93735 298072
rect 93596 298014 93735 298016
rect 94958 298014 95004 298074
rect 95068 298072 95115 298076
rect 95110 298016 95115 298072
rect 93596 298012 93602 298014
rect 93669 298011 93735 298014
rect 94998 298012 95004 298014
rect 95068 298012 95115 298016
rect 95049 298011 95115 298012
rect 82721 297938 82787 297941
rect 81758 297936 82787 297938
rect 81758 297880 82726 297936
rect 82782 297880 82787 297936
rect 81758 297878 82787 297880
rect 80348 297876 80354 297878
rect 81341 297875 81407 297878
rect 82721 297875 82787 297878
rect 83038 297876 83044 297940
rect 83108 297938 83114 297940
rect 84101 297938 84167 297941
rect 83108 297936 84167 297938
rect 83108 297880 84106 297936
rect 84162 297880 84167 297936
rect 83108 297878 84167 297880
rect 83108 297876 83114 297878
rect 84101 297875 84167 297878
rect 84510 297876 84516 297940
rect 84580 297938 84586 297940
rect 85389 297938 85455 297941
rect 84580 297936 85455 297938
rect 84580 297880 85394 297936
rect 85450 297880 85455 297936
rect 84580 297878 85455 297880
rect 84580 297876 84586 297878
rect 85389 297875 85455 297878
rect 86769 297938 86835 297941
rect 86902 297938 86908 297940
rect 86769 297936 86908 297938
rect 86769 297880 86774 297936
rect 86830 297880 86908 297936
rect 86769 297878 86908 297880
rect 86769 297875 86835 297878
rect 86902 297876 86908 297878
rect 86972 297876 86978 297940
rect 87638 297876 87644 297940
rect 87708 297938 87714 297940
rect 88241 297938 88307 297941
rect 87708 297936 88307 297938
rect 87708 297880 88246 297936
rect 88302 297880 88307 297936
rect 87708 297878 88307 297880
rect 87708 297876 87714 297878
rect 88241 297875 88307 297878
rect 90214 297876 90220 297940
rect 90284 297938 90290 297940
rect 90909 297938 90975 297941
rect 90284 297936 90975 297938
rect 90284 297880 90914 297936
rect 90970 297880 90975 297936
rect 90284 297878 90975 297880
rect 90284 297876 90290 297878
rect 90909 297875 90975 297878
rect 91318 297876 91324 297940
rect 91388 297938 91394 297940
rect 92381 297938 92447 297941
rect 91388 297936 92447 297938
rect 91388 297880 92386 297936
rect 92442 297880 92447 297936
rect 91388 297878 92447 297880
rect 91388 297876 91394 297878
rect 92381 297875 92447 297878
rect 93158 297876 93164 297940
rect 93228 297938 93234 297940
rect 93577 297938 93643 297941
rect 93228 297936 93643 297938
rect 93228 297880 93582 297936
rect 93638 297880 93643 297936
rect 93228 297878 93643 297880
rect 93228 297876 93234 297878
rect 93577 297875 93643 297878
rect 94446 297876 94452 297940
rect 94516 297938 94522 297940
rect 95141 297938 95207 297941
rect 94516 297936 95207 297938
rect 94516 297880 95146 297936
rect 95202 297880 95207 297936
rect 94516 297878 95207 297880
rect 95558 297938 95618 298148
rect 95926 298074 95986 298148
rect 96429 298074 96495 298077
rect 97073 298076 97139 298077
rect 97022 298074 97028 298076
rect 95926 298072 96495 298074
rect 95926 298016 96434 298072
rect 96490 298016 96495 298072
rect 95926 298014 96495 298016
rect 96982 298014 97028 298074
rect 97092 298072 97139 298076
rect 97134 298016 97139 298072
rect 96429 298011 96495 298014
rect 97022 298012 97028 298014
rect 97092 298012 97139 298016
rect 97073 298011 97139 298012
rect 97901 298076 97967 298077
rect 97901 298072 97948 298076
rect 98012 298074 98018 298076
rect 97901 298016 97906 298072
rect 97901 298012 97948 298016
rect 98012 298014 98058 298074
rect 98012 298012 98018 298014
rect 97901 298011 97967 298012
rect 96521 297938 96587 297941
rect 95558 297936 96587 297938
rect 95558 297880 96526 297936
rect 96582 297880 96587 297936
rect 95558 297878 96587 297880
rect 94516 297876 94522 297878
rect 95141 297875 95207 297878
rect 96521 297875 96587 297878
rect 96654 297876 96660 297940
rect 96724 297938 96730 297940
rect 97809 297938 97875 297941
rect 96724 297936 97875 297938
rect 96724 297880 97814 297936
rect 97870 297880 97875 297936
rect 96724 297878 97875 297880
rect 99422 297938 99482 298148
rect 102918 298077 102978 298148
rect 103286 298077 103346 298148
rect 100518 298012 100524 298076
rect 100588 298074 100594 298076
rect 100661 298074 100727 298077
rect 100588 298072 100727 298074
rect 100588 298016 100666 298072
rect 100722 298016 100727 298072
rect 100588 298014 100727 298016
rect 100588 298012 100594 298014
rect 100661 298011 100727 298014
rect 101438 298012 101444 298076
rect 101508 298074 101514 298076
rect 101857 298074 101923 298077
rect 101508 298072 101923 298074
rect 101508 298016 101862 298072
rect 101918 298016 101923 298072
rect 101508 298014 101923 298016
rect 102918 298072 103027 298077
rect 102918 298016 102966 298072
rect 103022 298016 103027 298072
rect 102918 298014 103027 298016
rect 103286 298072 103395 298077
rect 103286 298016 103334 298072
rect 103390 298016 103395 298072
rect 103286 298014 103395 298016
rect 101508 298012 101514 298014
rect 101857 298011 101923 298014
rect 102961 298011 103027 298014
rect 103329 298011 103395 298014
rect 104014 298012 104020 298076
rect 104084 298074 104090 298076
rect 104249 298074 104315 298077
rect 104084 298072 104315 298074
rect 104084 298016 104254 298072
rect 104310 298016 104315 298072
rect 104084 298014 104315 298016
rect 104084 298012 104090 298014
rect 104249 298011 104315 298014
rect 104382 298012 104388 298076
rect 104452 298074 104458 298076
rect 104709 298074 104775 298077
rect 104452 298072 104775 298074
rect 104452 298016 104714 298072
rect 104770 298016 104775 298072
rect 104452 298014 104775 298016
rect 104452 298012 104458 298014
rect 104709 298011 104775 298014
rect 105302 298012 105308 298076
rect 105372 298074 105378 298076
rect 105537 298074 105603 298077
rect 105372 298072 105603 298074
rect 105372 298016 105542 298072
rect 105598 298016 105603 298072
rect 105372 298014 105603 298016
rect 105372 298012 105378 298014
rect 105537 298011 105603 298014
rect 105670 298012 105676 298076
rect 105740 298074 105746 298076
rect 106089 298074 106155 298077
rect 106641 298076 106707 298077
rect 106590 298074 106596 298076
rect 105740 298072 106155 298074
rect 105740 298016 106094 298072
rect 106150 298016 106155 298072
rect 105740 298014 106155 298016
rect 106550 298014 106596 298074
rect 106660 298072 106707 298076
rect 106702 298016 106707 298072
rect 105740 298012 105746 298014
rect 106089 298011 106155 298014
rect 106590 298012 106596 298014
rect 106660 298012 106707 298016
rect 106958 298012 106964 298076
rect 107028 298074 107034 298076
rect 107469 298074 107535 298077
rect 107745 298076 107811 298077
rect 107694 298074 107700 298076
rect 107028 298072 107535 298074
rect 107028 298016 107474 298072
rect 107530 298016 107535 298072
rect 107028 298014 107535 298016
rect 107654 298014 107700 298074
rect 107764 298072 107811 298076
rect 107806 298016 107811 298072
rect 107028 298012 107034 298014
rect 106641 298011 106707 298012
rect 107469 298011 107535 298014
rect 107694 298012 107700 298014
rect 107764 298012 107811 298016
rect 107878 298012 107884 298076
rect 107948 298074 107954 298076
rect 108849 298074 108915 298077
rect 107948 298072 108915 298074
rect 107948 298016 108854 298072
rect 108910 298016 108915 298072
rect 107948 298014 108915 298016
rect 107948 298012 107954 298014
rect 107745 298011 107811 298012
rect 108849 298011 108915 298014
rect 109350 298012 109356 298076
rect 109420 298074 109426 298076
rect 110321 298074 110387 298077
rect 109420 298072 110387 298074
rect 109420 298016 110326 298072
rect 110382 298016 110387 298072
rect 109420 298014 110387 298016
rect 109420 298012 109426 298014
rect 110321 298011 110387 298014
rect 110638 298012 110644 298076
rect 110708 298074 110714 298076
rect 111609 298074 111675 298077
rect 110708 298072 111675 298074
rect 110708 298016 111614 298072
rect 111670 298016 111675 298072
rect 110708 298014 111675 298016
rect 110708 298012 110714 298014
rect 111609 298011 111675 298014
rect 112989 298076 113055 298077
rect 112989 298072 113036 298076
rect 113100 298074 113106 298076
rect 112989 298016 112994 298072
rect 112989 298012 113036 298016
rect 113100 298014 113146 298074
rect 113100 298012 113106 298014
rect 114318 298012 114324 298076
rect 114388 298074 114394 298076
rect 114461 298074 114527 298077
rect 114388 298072 114527 298074
rect 114388 298016 114466 298072
rect 114522 298016 114527 298072
rect 114388 298014 114527 298016
rect 114388 298012 114394 298014
rect 112989 298011 113055 298012
rect 114461 298011 114527 298014
rect 115606 298012 115612 298076
rect 115676 298074 115682 298076
rect 115841 298074 115907 298077
rect 115676 298072 115907 298074
rect 115676 298016 115846 298072
rect 115902 298016 115907 298072
rect 115676 298014 115907 298016
rect 115676 298012 115682 298014
rect 115841 298011 115907 298014
rect 116894 298012 116900 298076
rect 116964 298074 116970 298076
rect 117221 298074 117287 298077
rect 116964 298072 117287 298074
rect 116964 298016 117226 298072
rect 117282 298016 117287 298072
rect 116964 298014 117287 298016
rect 116964 298012 116970 298014
rect 117221 298011 117287 298014
rect 215845 298076 215911 298077
rect 215845 298072 215892 298076
rect 215956 298074 215962 298076
rect 224953 298074 225019 298077
rect 225462 298074 225522 298148
rect 257846 298077 257906 298148
rect 215845 298016 215850 298072
rect 215845 298012 215892 298016
rect 215956 298014 216002 298074
rect 224953 298072 225522 298074
rect 224953 298016 224958 298072
rect 225014 298016 225522 298072
rect 224953 298014 225522 298016
rect 226333 298074 226399 298077
rect 226742 298074 226748 298076
rect 226333 298072 226748 298074
rect 226333 298016 226338 298072
rect 226394 298016 226748 298072
rect 226333 298014 226748 298016
rect 215956 298012 215962 298014
rect 215845 298011 215911 298012
rect 224953 298011 225019 298014
rect 226333 298011 226399 298014
rect 226742 298012 226748 298014
rect 226812 298012 226818 298076
rect 227713 298074 227779 298077
rect 227846 298074 227852 298076
rect 227713 298072 227852 298074
rect 227713 298016 227718 298072
rect 227774 298016 227852 298072
rect 227713 298014 227852 298016
rect 227713 298011 227779 298014
rect 227846 298012 227852 298014
rect 227916 298012 227922 298076
rect 230473 298074 230539 298077
rect 231342 298074 231348 298076
rect 230473 298072 231348 298074
rect 230473 298016 230478 298072
rect 230534 298016 231348 298072
rect 230473 298014 231348 298016
rect 230473 298011 230539 298014
rect 231342 298012 231348 298014
rect 231412 298012 231418 298076
rect 231945 298074 232011 298077
rect 232630 298074 232636 298076
rect 231945 298072 232636 298074
rect 231945 298016 231950 298072
rect 232006 298016 232636 298072
rect 231945 298014 232636 298016
rect 231945 298011 232011 298014
rect 232630 298012 232636 298014
rect 232700 298012 232706 298076
rect 233233 298074 233299 298077
rect 233550 298074 233556 298076
rect 233233 298072 233556 298074
rect 233233 298016 233238 298072
rect 233294 298016 233556 298072
rect 233233 298014 233556 298016
rect 233233 298011 233299 298014
rect 233550 298012 233556 298014
rect 233620 298012 233626 298076
rect 234705 298074 234771 298077
rect 237189 298076 237255 298077
rect 235022 298074 235028 298076
rect 234705 298072 235028 298074
rect 234705 298016 234710 298072
rect 234766 298016 235028 298072
rect 234705 298014 235028 298016
rect 234705 298011 234771 298014
rect 235022 298012 235028 298014
rect 235092 298012 235098 298076
rect 237189 298072 237236 298076
rect 237300 298074 237306 298076
rect 237189 298016 237194 298072
rect 237189 298012 237236 298016
rect 237300 298014 237346 298074
rect 237300 298012 237306 298014
rect 238334 298012 238340 298076
rect 238404 298074 238410 298076
rect 238661 298074 238727 298077
rect 238404 298072 238727 298074
rect 238404 298016 238666 298072
rect 238722 298016 238727 298072
rect 238404 298014 238727 298016
rect 238404 298012 238410 298014
rect 237189 298011 237255 298012
rect 238661 298011 238727 298014
rect 240133 298074 240199 298077
rect 240358 298074 240364 298076
rect 240133 298072 240364 298074
rect 240133 298016 240138 298072
rect 240194 298016 240364 298072
rect 240133 298014 240364 298016
rect 240133 298011 240199 298014
rect 240358 298012 240364 298014
rect 240428 298012 240434 298076
rect 240726 298012 240732 298076
rect 240796 298074 240802 298076
rect 241421 298074 241487 298077
rect 240796 298072 241487 298074
rect 240796 298016 241426 298072
rect 241482 298016 241487 298072
rect 240796 298014 241487 298016
rect 240796 298012 240802 298014
rect 241421 298011 241487 298014
rect 242893 298076 242959 298077
rect 244089 298076 244155 298077
rect 242893 298072 242940 298076
rect 243004 298074 243010 298076
rect 244038 298074 244044 298076
rect 242893 298016 242898 298072
rect 242893 298012 242940 298016
rect 243004 298014 243050 298074
rect 243998 298014 244044 298074
rect 244108 298072 244155 298076
rect 244150 298016 244155 298072
rect 243004 298012 243010 298014
rect 244038 298012 244044 298014
rect 244108 298012 244155 298016
rect 242893 298011 242959 298012
rect 244089 298011 244155 298012
rect 244273 298074 244339 298077
rect 245561 298076 245627 298077
rect 246849 298076 246915 298077
rect 244406 298074 244412 298076
rect 244273 298072 244412 298074
rect 244273 298016 244278 298072
rect 244334 298016 244412 298072
rect 244273 298014 244412 298016
rect 244273 298011 244339 298014
rect 244406 298012 244412 298014
rect 244476 298012 244482 298076
rect 245510 298074 245516 298076
rect 245470 298014 245516 298074
rect 245580 298072 245627 298076
rect 246798 298074 246804 298076
rect 245622 298016 245627 298072
rect 245510 298012 245516 298014
rect 245580 298012 245627 298016
rect 246758 298014 246804 298074
rect 246868 298072 246915 298076
rect 246910 298016 246915 298072
rect 246798 298012 246804 298014
rect 246868 298012 246915 298016
rect 247902 298012 247908 298076
rect 247972 298074 247978 298076
rect 248229 298074 248295 298077
rect 247972 298072 248295 298074
rect 247972 298016 248234 298072
rect 248290 298016 248295 298072
rect 247972 298014 248295 298016
rect 247972 298012 247978 298014
rect 245561 298011 245627 298012
rect 246849 298011 246915 298012
rect 248229 298011 248295 298014
rect 249374 298012 249380 298076
rect 249444 298074 249450 298076
rect 249701 298074 249767 298077
rect 249444 298072 249767 298074
rect 249444 298016 249706 298072
rect 249762 298016 249767 298072
rect 249444 298014 249767 298016
rect 249444 298012 249450 298014
rect 249701 298011 249767 298014
rect 250662 298012 250668 298076
rect 250732 298074 250738 298076
rect 250989 298074 251055 298077
rect 250732 298072 251055 298074
rect 250732 298016 250994 298072
rect 251050 298016 251055 298072
rect 250732 298014 251055 298016
rect 250732 298012 250738 298014
rect 250989 298011 251055 298014
rect 252369 298074 252435 298077
rect 252502 298074 252508 298076
rect 252369 298072 252508 298074
rect 252369 298016 252374 298072
rect 252430 298016 252508 298072
rect 252369 298014 252508 298016
rect 252369 298011 252435 298014
rect 252502 298012 252508 298014
rect 252572 298012 252578 298076
rect 253606 298012 253612 298076
rect 253676 298074 253682 298076
rect 253749 298074 253815 298077
rect 253676 298072 253815 298074
rect 253676 298016 253754 298072
rect 253810 298016 253815 298072
rect 253676 298014 253815 298016
rect 253676 298012 253682 298014
rect 253749 298011 253815 298014
rect 254894 298012 254900 298076
rect 254964 298074 254970 298076
rect 255129 298074 255195 298077
rect 254964 298072 255195 298074
rect 254964 298016 255134 298072
rect 255190 298016 255195 298072
rect 254964 298014 255195 298016
rect 254964 298012 254970 298014
rect 255129 298011 255195 298014
rect 255998 298012 256004 298076
rect 256068 298074 256074 298076
rect 256509 298074 256575 298077
rect 256068 298072 256575 298074
rect 256068 298016 256514 298072
rect 256570 298016 256575 298072
rect 256068 298014 256575 298016
rect 257846 298072 257955 298077
rect 257846 298016 257894 298072
rect 257950 298016 257955 298072
rect 257846 298014 257955 298016
rect 256068 298012 256074 298014
rect 256509 298011 256575 298014
rect 257889 298011 257955 298014
rect 259177 298074 259243 298077
rect 259310 298074 259316 298076
rect 259177 298072 259316 298074
rect 259177 298016 259182 298072
rect 259238 298016 259316 298072
rect 259177 298014 259316 298016
rect 259177 298011 259243 298014
rect 259310 298012 259316 298014
rect 259380 298012 259386 298076
rect 260649 298074 260715 298077
rect 260782 298074 260788 298076
rect 260649 298072 260788 298074
rect 260649 298016 260654 298072
rect 260710 298016 260788 298072
rect 260649 298014 260788 298016
rect 260649 298011 260715 298014
rect 260782 298012 260788 298014
rect 260852 298012 260858 298076
rect 100569 297938 100635 297941
rect 99422 297936 100635 297938
rect 99422 297880 100574 297936
rect 100630 297880 100635 297936
rect 99422 297878 100635 297880
rect 96724 297876 96730 297878
rect 97809 297875 97875 297878
rect 100569 297875 100635 297878
rect 100702 297876 100708 297940
rect 100772 297938 100778 297940
rect 101949 297938 102015 297941
rect 100772 297936 102015 297938
rect 100772 297880 101954 297936
rect 102010 297880 102015 297936
rect 100772 297878 102015 297880
rect 100772 297876 100778 297878
rect 101949 297875 102015 297878
rect 111926 297876 111932 297940
rect 111996 297938 112002 297940
rect 113081 297938 113147 297941
rect 111996 297936 113147 297938
rect 111996 297880 113086 297936
rect 113142 297880 113147 297936
rect 111996 297878 113147 297880
rect 111996 297876 112002 297878
rect 113081 297875 113147 297878
rect 237373 297938 237439 297941
rect 237782 297938 237788 297940
rect 237373 297936 237788 297938
rect 237373 297880 237378 297936
rect 237434 297880 237788 297936
rect 237373 297878 237788 297880
rect 237373 297875 237439 297878
rect 237782 297876 237788 297878
rect 237852 297876 237858 297940
rect 238753 297938 238819 297941
rect 239254 297938 239260 297940
rect 238753 297936 239260 297938
rect 238753 297880 238758 297936
rect 238814 297880 239260 297936
rect 238753 297878 239260 297880
rect 238753 297875 238819 297878
rect 239254 297876 239260 297878
rect 239324 297876 239330 297940
rect 241513 297938 241579 297941
rect 242014 297938 242020 297940
rect 241513 297936 242020 297938
rect 241513 297880 241518 297936
rect 241574 297880 242020 297936
rect 241513 297878 242020 297880
rect 241513 297875 241579 297878
rect 242014 297876 242020 297878
rect 242084 297876 242090 297940
rect 243077 297938 243143 297941
rect 244181 297938 244247 297941
rect 243077 297936 244247 297938
rect 243077 297880 243082 297936
rect 243138 297880 244186 297936
rect 244242 297880 244247 297936
rect 243077 297878 244247 297880
rect 243077 297875 243143 297878
rect 244181 297875 244247 297878
rect 245694 297876 245700 297940
rect 245764 297938 245770 297940
rect 246757 297938 246823 297941
rect 245764 297936 246823 297938
rect 245764 297880 246762 297936
rect 246818 297880 246823 297936
rect 245764 297878 246823 297880
rect 245764 297876 245770 297878
rect 246757 297875 246823 297878
rect 247718 297876 247724 297940
rect 247788 297938 247794 297940
rect 248321 297938 248387 297941
rect 247788 297936 248387 297938
rect 247788 297880 248326 297936
rect 248382 297880 248387 297936
rect 247788 297878 248387 297880
rect 247788 297876 247794 297878
rect 248321 297875 248387 297878
rect 249006 297876 249012 297940
rect 249076 297938 249082 297940
rect 249609 297938 249675 297941
rect 249076 297936 249675 297938
rect 249076 297880 249614 297936
rect 249670 297880 249675 297936
rect 249076 297878 249675 297880
rect 249076 297876 249082 297878
rect 249609 297875 249675 297878
rect 250294 297876 250300 297940
rect 250364 297938 250370 297940
rect 251081 297938 251147 297941
rect 250364 297936 251147 297938
rect 250364 297880 251086 297936
rect 251142 297880 251147 297936
rect 250364 297878 251147 297880
rect 250364 297876 250370 297878
rect 251081 297875 251147 297878
rect 251398 297876 251404 297940
rect 251468 297938 251474 297940
rect 252277 297938 252343 297941
rect 251468 297936 252343 297938
rect 251468 297880 252282 297936
rect 252338 297880 252343 297936
rect 251468 297878 252343 297880
rect 251468 297876 251474 297878
rect 252277 297875 252343 297878
rect 253054 297876 253060 297940
rect 253124 297938 253130 297940
rect 253841 297938 253907 297941
rect 253124 297936 253907 297938
rect 253124 297880 253846 297936
rect 253902 297880 253907 297936
rect 253124 297878 253907 297880
rect 253124 297876 253130 297878
rect 253841 297875 253907 297878
rect 254526 297876 254532 297940
rect 254596 297938 254602 297940
rect 255221 297938 255287 297941
rect 254596 297936 255287 297938
rect 254596 297880 255226 297936
rect 255282 297880 255287 297936
rect 254596 297878 255287 297880
rect 254596 297876 254602 297878
rect 255221 297875 255287 297878
rect 255630 297876 255636 297940
rect 255700 297938 255706 297940
rect 256601 297938 256667 297941
rect 255700 297936 256667 297938
rect 255700 297880 256606 297936
rect 256662 297880 256667 297936
rect 255700 297878 256667 297880
rect 255700 297876 255706 297878
rect 256601 297875 256667 297878
rect 257102 297876 257108 297940
rect 257172 297938 257178 297940
rect 257797 297938 257863 297941
rect 257172 297936 257863 297938
rect 257172 297880 257802 297936
rect 257858 297880 257863 297936
rect 257172 297878 257863 297880
rect 257172 297876 257178 297878
rect 257797 297875 257863 297878
rect 259126 297876 259132 297940
rect 259196 297938 259202 297940
rect 259361 297938 259427 297941
rect 259196 297936 259427 297938
rect 259196 297880 259366 297936
rect 259422 297880 259427 297936
rect 259196 297878 259427 297880
rect 259196 297876 259202 297878
rect 259361 297875 259427 297878
rect 260598 297876 260604 297940
rect 260668 297938 260674 297940
rect 260741 297938 260807 297941
rect 260668 297936 260807 297938
rect 260668 297880 260746 297936
rect 260802 297880 260807 297936
rect 260668 297878 260807 297880
rect 261526 297938 261586 298148
rect 261894 298074 261954 298148
rect 262029 298074 262095 298077
rect 261894 298072 262095 298074
rect 261894 298016 262034 298072
rect 262090 298016 262095 298072
rect 261894 298014 262095 298016
rect 262029 298011 262095 298014
rect 263174 298012 263180 298076
rect 263244 298074 263250 298076
rect 263501 298074 263567 298077
rect 263244 298072 263567 298074
rect 263244 298016 263506 298072
rect 263562 298016 263567 298072
rect 263244 298014 263567 298016
rect 265206 298074 265266 298148
rect 266169 298074 266235 298077
rect 265206 298072 266235 298074
rect 265206 298016 266174 298072
rect 266230 298016 266235 298072
rect 265206 298014 266235 298016
rect 271830 298074 271890 298148
rect 273069 298074 273135 298077
rect 271830 298072 273135 298074
rect 271830 298016 273074 298072
rect 273130 298016 273135 298072
rect 271830 298014 273135 298016
rect 263244 298012 263250 298014
rect 263501 298011 263567 298014
rect 266169 298011 266235 298014
rect 273069 298011 273135 298014
rect 274398 298012 274404 298076
rect 274468 298074 274474 298076
rect 274541 298074 274607 298077
rect 274468 298072 274607 298074
rect 274468 298016 274546 298072
rect 274602 298016 274607 298072
rect 274468 298014 274607 298016
rect 275510 298074 275570 298148
rect 275921 298074 275987 298077
rect 275510 298072 275987 298074
rect 275510 298016 275926 298072
rect 275982 298016 275987 298072
rect 275510 298014 275987 298016
rect 274468 298012 274474 298014
rect 274541 298011 274607 298014
rect 275921 298011 275987 298014
rect 276790 298012 276796 298076
rect 276860 298074 276866 298076
rect 277301 298074 277367 298077
rect 276860 298072 277367 298074
rect 276860 298016 277306 298072
rect 277362 298016 277367 298072
rect 276860 298014 277367 298016
rect 276860 298012 276866 298014
rect 277301 298011 277367 298014
rect 262121 297938 262187 297941
rect 261526 297936 262187 297938
rect 261526 297880 262126 297936
rect 262182 297880 262187 297936
rect 261526 297878 262187 297880
rect 260668 297876 260674 297878
rect 260741 297875 260807 297878
rect 262121 297875 262187 297878
rect 262990 297876 262996 297940
rect 263060 297938 263066 297940
rect 263409 297938 263475 297941
rect 263060 297936 263475 297938
rect 263060 297880 263414 297936
rect 263470 297880 263475 297936
rect 263060 297878 263475 297880
rect 263060 297876 263066 297878
rect 263409 297875 263475 297878
rect 85798 297740 85804 297804
rect 85868 297802 85874 297804
rect 86861 297802 86927 297805
rect 85868 297800 86927 297802
rect 85868 297744 86866 297800
rect 86922 297744 86927 297800
rect 85868 297742 86927 297744
rect 85868 297740 85874 297742
rect 86861 297739 86927 297742
rect 92606 297740 92612 297804
rect 92676 297802 92682 297804
rect 93761 297802 93827 297805
rect 92676 297800 93827 297802
rect 92676 297744 93766 297800
rect 93822 297744 93827 297800
rect 92676 297742 93827 297744
rect 92676 297740 92682 297742
rect 93761 297739 93827 297742
rect 101806 297740 101812 297804
rect 101876 297802 101882 297804
rect 102041 297802 102107 297805
rect 101876 297800 102107 297802
rect 101876 297744 102046 297800
rect 102102 297744 102107 297800
rect 101876 297742 102107 297744
rect 101876 297740 101882 297742
rect 102041 297739 102107 297742
rect 229277 297802 229343 297805
rect 230054 297802 230060 297804
rect 229277 297800 230060 297802
rect 229277 297744 229282 297800
rect 229338 297744 230060 297800
rect 229277 297742 230060 297744
rect 229277 297739 229343 297742
rect 230054 297740 230060 297742
rect 230124 297740 230130 297804
rect 236494 297740 236500 297804
rect 236564 297802 236570 297804
rect 237281 297802 237347 297805
rect 236564 297800 237347 297802
rect 236564 297744 237286 297800
rect 237342 297744 237347 297800
rect 236564 297742 237347 297744
rect 236564 297740 236570 297742
rect 237281 297739 237347 297742
rect 241830 297740 241836 297804
rect 241900 297802 241906 297804
rect 242801 297802 242867 297805
rect 241900 297800 242867 297802
rect 241900 297744 242806 297800
rect 242862 297744 242867 297800
rect 241900 297742 242867 297744
rect 241900 297740 241906 297742
rect 242801 297739 242867 297742
rect 246614 297740 246620 297804
rect 246684 297802 246690 297804
rect 246941 297802 247007 297805
rect 246684 297800 247007 297802
rect 246684 297744 246946 297800
rect 247002 297744 247007 297800
rect 246684 297742 247007 297744
rect 246684 297740 246690 297742
rect 246941 297739 247007 297742
rect 251950 297740 251956 297804
rect 252020 297802 252026 297804
rect 252461 297802 252527 297805
rect 252020 297800 252527 297802
rect 252020 297744 252466 297800
rect 252522 297744 252527 297800
rect 252020 297742 252527 297744
rect 252020 297740 252026 297742
rect 252461 297739 252527 297742
rect 256734 297740 256740 297804
rect 256804 297802 256810 297804
rect 257981 297802 258047 297805
rect 256804 297800 258047 297802
rect 256804 297744 257986 297800
rect 258042 297744 258047 297800
rect 256804 297742 258047 297744
rect 256804 297740 256810 297742
rect 257981 297739 258047 297742
rect 258390 297740 258396 297804
rect 258460 297802 258466 297804
rect 259269 297802 259335 297805
rect 258460 297800 259335 297802
rect 258460 297744 259274 297800
rect 259330 297744 259335 297800
rect 258460 297742 259335 297744
rect 258460 297740 258466 297742
rect 259269 297739 259335 297742
rect 99046 297468 99052 297532
rect 99116 297530 99122 297532
rect 408534 297530 408540 297532
rect 99116 297470 408540 297530
rect 99116 297468 99122 297470
rect 408534 297468 408540 297470
rect 408604 297468 408610 297532
rect 98310 297332 98316 297396
rect 98380 297394 98386 297396
rect 408718 297394 408724 297396
rect 98380 297334 408724 297394
rect 98380 297332 98386 297334
rect 408718 297332 408724 297334
rect 408788 297332 408794 297396
rect 83958 297060 83964 297124
rect 84028 297122 84034 297124
rect 85297 297122 85363 297125
rect 84028 297120 85363 297122
rect 84028 297064 85302 297120
rect 85358 297064 85363 297120
rect 84028 297062 85363 297064
rect 84028 297060 84034 297062
rect 85297 297059 85363 297062
rect 238569 297122 238635 297125
rect 240041 297122 240107 297125
rect 238569 297120 240107 297122
rect 238569 297064 238574 297120
rect 238630 297064 240046 297120
rect 240102 297064 240107 297120
rect 238569 297062 240107 297064
rect 238569 297059 238635 297062
rect 240041 297059 240107 297062
rect 266854 297060 266860 297124
rect 266924 297122 266930 297124
rect 267641 297122 267707 297125
rect 266924 297120 267707 297122
rect 266924 297064 267646 297120
rect 267702 297064 267707 297120
rect 266924 297062 267707 297064
rect 266924 297060 266930 297062
rect 267641 297059 267707 297062
rect 264094 296924 264100 296988
rect 264164 296986 264170 296988
rect 264789 296986 264855 296989
rect 264164 296984 264855 296986
rect 264164 296928 264794 296984
rect 264850 296928 264855 296984
rect 264164 296926 264855 296928
rect 264164 296924 264170 296926
rect 264789 296923 264855 296926
rect 266670 296924 266676 296988
rect 266740 296986 266746 296988
rect 267457 296986 267523 296989
rect 266740 296984 267523 296986
rect 266740 296928 267462 296984
rect 267518 296928 267523 296984
rect 266740 296926 267523 296928
rect 266740 296924 266746 296926
rect 267457 296923 267523 296926
rect 264462 296788 264468 296852
rect 264532 296850 264538 296852
rect 264881 296850 264947 296853
rect 264532 296848 264947 296850
rect 264532 296792 264886 296848
rect 264942 296792 264947 296848
rect 264532 296790 264947 296792
rect 264532 296788 264538 296790
rect 264881 296787 264947 296790
rect 265750 296788 265756 296852
rect 265820 296850 265826 296852
rect 266261 296850 266327 296853
rect 267549 296852 267615 296853
rect 267549 296850 267596 296852
rect 265820 296848 266327 296850
rect 265820 296792 266266 296848
rect 266322 296792 266327 296848
rect 265820 296790 266327 296792
rect 267504 296848 267596 296850
rect 267504 296792 267554 296848
rect 267504 296790 267596 296792
rect 265820 296788 265826 296790
rect 266261 296787 266327 296790
rect 267549 296788 267596 296790
rect 267660 296788 267666 296852
rect 267958 296788 267964 296852
rect 268028 296850 268034 296852
rect 269021 296850 269087 296853
rect 268028 296848 269087 296850
rect 268028 296792 269026 296848
rect 269082 296792 269087 296848
rect 268028 296790 269087 296792
rect 268028 296788 268034 296790
rect 267549 296787 267615 296788
rect 269021 296787 269087 296790
rect 269246 296788 269252 296852
rect 269316 296850 269322 296852
rect 270401 296850 270467 296853
rect 269316 296848 270467 296850
rect 269316 296792 270406 296848
rect 270462 296792 270467 296848
rect 269316 296790 270467 296792
rect 269316 296788 269322 296790
rect 270401 296787 270467 296790
rect 270534 296788 270540 296852
rect 270604 296850 270610 296852
rect 271781 296850 271847 296853
rect 273161 296852 273227 296853
rect 273110 296850 273116 296852
rect 270604 296848 271847 296850
rect 270604 296792 271786 296848
rect 271842 296792 271847 296848
rect 270604 296790 271847 296792
rect 273070 296790 273116 296850
rect 273180 296848 273227 296852
rect 273222 296792 273227 296848
rect 270604 296788 270610 296790
rect 271781 296787 271847 296790
rect 273110 296788 273116 296790
rect 273180 296788 273227 296792
rect 273161 296787 273227 296788
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 408953 251834 409019 251837
rect 409270 251834 409276 251836
rect 408953 251832 409276 251834
rect 408953 251776 408958 251832
rect 409014 251776 409276 251832
rect 408953 251774 409276 251776
rect 408953 251771 409019 251774
rect 409270 251772 409276 251774
rect 409340 251772 409346 251836
rect 408861 249658 408927 249661
rect 408861 249656 409338 249658
rect 408861 249600 408866 249656
rect 408922 249600 409338 249656
rect 408861 249598 409338 249600
rect 408861 249595 408927 249598
rect 186313 249522 186379 249525
rect 186313 249520 190164 249522
rect 186313 249464 186318 249520
rect 186374 249464 190164 249520
rect 186313 249462 190164 249464
rect 186313 249459 186379 249462
rect 409278 249084 409338 249598
rect 186313 248298 186379 248301
rect 186313 248296 190164 248298
rect 186313 248240 186318 248296
rect 186374 248240 190164 248296
rect 186313 248238 190164 248240
rect 186313 248235 186379 248238
rect 409270 248236 409276 248300
rect 409340 248298 409346 248300
rect 409413 248298 409479 248301
rect 409340 248296 409479 248298
rect 409340 248240 409418 248296
rect 409474 248240 409479 248296
rect 409340 248238 409479 248240
rect 409340 248236 409346 248238
rect 409413 248235 409479 248238
rect 409321 247754 409387 247757
rect 409321 247752 409522 247754
rect 409321 247696 409326 247752
rect 409382 247696 409522 247752
rect 409321 247694 409522 247696
rect 409321 247691 409387 247694
rect 186405 247210 186471 247213
rect 186405 247208 190164 247210
rect 186405 247152 186410 247208
rect 186466 247152 190164 247208
rect 409462 247180 409522 247694
rect 186405 247150 190164 247152
rect 186405 247147 186471 247150
rect 186313 245986 186379 245989
rect 186313 245984 190164 245986
rect 186313 245928 186318 245984
rect 186374 245928 190164 245984
rect 186313 245926 190164 245928
rect 186313 245923 186379 245926
rect 409321 245578 409387 245581
rect 409278 245576 409387 245578
rect 409278 245520 409326 245576
rect 409382 245520 409387 245576
rect 409278 245515 409387 245520
rect 409278 245276 409338 245515
rect 583520 245428 584960 245668
rect 186313 244898 186379 244901
rect 186313 244896 190164 244898
rect 186313 244840 186318 244896
rect 186374 244840 190164 244896
rect 186313 244838 190164 244840
rect 186313 244835 186379 244838
rect 186313 243674 186379 243677
rect 409321 243674 409387 243677
rect 186313 243672 190164 243674
rect 186313 243616 186318 243672
rect 186374 243616 190164 243672
rect 186313 243614 190164 243616
rect 409278 243672 409387 243674
rect 409278 243616 409326 243672
rect 409382 243616 409387 243672
rect 186313 243611 186379 243614
rect 409278 243611 409387 243616
rect 409278 243372 409338 243611
rect 186313 242586 186379 242589
rect 186313 242584 190164 242586
rect 186313 242528 186318 242584
rect 186374 242528 190164 242584
rect 186313 242526 190164 242528
rect 186313 242523 186379 242526
rect 409321 241634 409387 241637
rect 409321 241632 409522 241634
rect 409321 241576 409326 241632
rect 409382 241576 409522 241632
rect 409321 241574 409522 241576
rect 409321 241571 409387 241574
rect 409462 241468 409522 241574
rect 186313 241362 186379 241365
rect 186313 241360 190164 241362
rect 186313 241304 186318 241360
rect 186374 241304 190164 241360
rect 186313 241302 190164 241304
rect 186313 241299 186379 241302
rect -960 240940 480 241180
rect 186313 240138 186379 240141
rect 186313 240136 190164 240138
rect 186313 240080 186318 240136
rect 186374 240080 190164 240136
rect 186313 240078 190164 240080
rect 186313 240075 186379 240078
rect 410517 239594 410583 239597
rect 409860 239592 410583 239594
rect 409860 239536 410522 239592
rect 410578 239536 410583 239592
rect 409860 239534 410583 239536
rect 410517 239531 410583 239534
rect 186405 239050 186471 239053
rect 186405 239048 190164 239050
rect 186405 238992 186410 239048
rect 186466 238992 190164 239048
rect 186405 238990 190164 238992
rect 186405 238987 186471 238990
rect 187141 237826 187207 237829
rect 187141 237824 190164 237826
rect 187141 237768 187146 237824
rect 187202 237768 190164 237824
rect 187141 237766 190164 237768
rect 187141 237763 187207 237766
rect 409270 237764 409276 237828
rect 409340 237826 409346 237828
rect 409340 237766 409522 237826
rect 409340 237764 409346 237766
rect 409462 237660 409522 237766
rect 186313 236738 186379 236741
rect 186313 236736 190164 236738
rect 186313 236680 186318 236736
rect 186374 236680 190164 236736
rect 186313 236678 190164 236680
rect 186313 236675 186379 236678
rect 411897 235786 411963 235789
rect 409860 235784 411963 235786
rect 409860 235728 411902 235784
rect 411958 235728 411963 235784
rect 409860 235726 411963 235728
rect 411897 235723 411963 235726
rect 186313 235514 186379 235517
rect 186313 235512 190164 235514
rect 186313 235456 186318 235512
rect 186374 235456 190164 235512
rect 186313 235454 190164 235456
rect 186313 235451 186379 235454
rect 186313 234426 186379 234429
rect 186313 234424 190164 234426
rect 186313 234368 186318 234424
rect 186374 234368 190164 234424
rect 186313 234366 190164 234368
rect 186313 234363 186379 234366
rect 409270 234228 409276 234292
rect 409340 234228 409346 234292
rect 409278 233852 409338 234228
rect 186313 233202 186379 233205
rect 186313 233200 190164 233202
rect 186313 233144 186318 233200
rect 186374 233144 190164 233200
rect 186313 233142 190164 233144
rect 186313 233139 186379 233142
rect 583520 232236 584960 232476
rect 186405 232114 186471 232117
rect 186405 232112 190164 232114
rect 186405 232056 186410 232112
rect 186466 232056 190164 232112
rect 186405 232054 190164 232056
rect 186405 232051 186471 232054
rect 410425 231978 410491 231981
rect 409860 231976 410491 231978
rect 409860 231920 410430 231976
rect 410486 231920 410491 231976
rect 409860 231918 410491 231920
rect 410425 231915 410491 231918
rect 186313 230890 186379 230893
rect 186313 230888 190164 230890
rect 186313 230832 186318 230888
rect 186374 230832 190164 230888
rect 186313 230830 190164 230832
rect 186313 230827 186379 230830
rect 411621 230074 411687 230077
rect 409860 230072 411687 230074
rect 409860 230016 411626 230072
rect 411682 230016 411687 230072
rect 409860 230014 411687 230016
rect 411621 230011 411687 230014
rect 186313 229666 186379 229669
rect 186313 229664 190164 229666
rect 186313 229608 186318 229664
rect 186374 229608 190164 229664
rect 186313 229606 190164 229608
rect 186313 229603 186379 229606
rect 186313 228578 186379 228581
rect 186313 228576 190164 228578
rect 186313 228520 186318 228576
rect 186374 228520 190164 228576
rect 186313 228518 190164 228520
rect 186313 228515 186379 228518
rect 410241 228170 410307 228173
rect 409860 228168 410307 228170
rect -960 227884 480 228124
rect 409860 228112 410246 228168
rect 410302 228112 410307 228168
rect 409860 228110 410307 228112
rect 410241 228107 410307 228110
rect 186313 227354 186379 227357
rect 186313 227352 190164 227354
rect 186313 227296 186318 227352
rect 186374 227296 190164 227352
rect 186313 227294 190164 227296
rect 186313 227291 186379 227294
rect 186405 226266 186471 226269
rect 410333 226266 410399 226269
rect 186405 226264 190164 226266
rect 186405 226208 186410 226264
rect 186466 226208 190164 226264
rect 186405 226206 190164 226208
rect 409860 226264 410399 226266
rect 409860 226208 410338 226264
rect 410394 226208 410399 226264
rect 409860 226206 410399 226208
rect 186405 226203 186471 226206
rect 410333 226203 410399 226206
rect 186313 225042 186379 225045
rect 186313 225040 190164 225042
rect 186313 224984 186318 225040
rect 186374 224984 190164 225040
rect 186313 224982 190164 224984
rect 186313 224979 186379 224982
rect 410149 224362 410215 224365
rect 409860 224360 410215 224362
rect 409860 224304 410154 224360
rect 410210 224304 410215 224360
rect 409860 224302 410215 224304
rect 410149 224299 410215 224302
rect 186313 223954 186379 223957
rect 186313 223952 190164 223954
rect 186313 223896 186318 223952
rect 186374 223896 190164 223952
rect 186313 223894 190164 223896
rect 186313 223891 186379 223894
rect 186313 222730 186379 222733
rect 186313 222728 190164 222730
rect 186313 222672 186318 222728
rect 186374 222672 190164 222728
rect 186313 222670 190164 222672
rect 186313 222667 186379 222670
rect 411805 222458 411871 222461
rect 409860 222456 411871 222458
rect 409860 222400 411810 222456
rect 411866 222400 411871 222456
rect 409860 222398 411871 222400
rect 411805 222395 411871 222398
rect 186313 221506 186379 221509
rect 186313 221504 190164 221506
rect 186313 221448 186318 221504
rect 186374 221448 190164 221504
rect 186313 221446 190164 221448
rect 186313 221443 186379 221446
rect 411529 220554 411595 220557
rect 409860 220552 411595 220554
rect 409860 220496 411534 220552
rect 411590 220496 411595 220552
rect 409860 220494 411595 220496
rect 411529 220491 411595 220494
rect 186313 220418 186379 220421
rect 186313 220416 190164 220418
rect 186313 220360 186318 220416
rect 186374 220360 190164 220416
rect 186313 220358 190164 220360
rect 186313 220355 186379 220358
rect 186405 219194 186471 219197
rect 186405 219192 190164 219194
rect 186405 219136 186410 219192
rect 186466 219136 190164 219192
rect 186405 219134 190164 219136
rect 186405 219131 186471 219134
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 411713 218650 411779 218653
rect 409860 218648 411779 218650
rect 409860 218592 411718 218648
rect 411774 218592 411779 218648
rect 409860 218590 411779 218592
rect 411713 218587 411779 218590
rect 186313 218106 186379 218109
rect 186313 218104 190164 218106
rect 186313 218048 186318 218104
rect 186374 218048 190164 218104
rect 186313 218046 190164 218048
rect 186313 218043 186379 218046
rect 409965 217290 410031 217293
rect 409830 217288 410031 217290
rect 409830 217232 409970 217288
rect 410026 217232 410031 217288
rect 409830 217230 410031 217232
rect 186313 216882 186379 216885
rect 186313 216880 190164 216882
rect 186313 216824 186318 216880
rect 186374 216824 190164 216880
rect 186313 216822 190164 216824
rect 186313 216819 186379 216822
rect 409830 216716 409890 217230
rect 409965 217227 410031 217230
rect 186313 215794 186379 215797
rect 186313 215792 190164 215794
rect 186313 215736 186318 215792
rect 186374 215736 190164 215792
rect 186313 215734 190164 215736
rect 186313 215731 186379 215734
rect -960 214828 480 215068
rect 411345 214842 411411 214845
rect 409860 214840 411411 214842
rect 409860 214784 411350 214840
rect 411406 214784 411411 214840
rect 409860 214782 411411 214784
rect 411345 214779 411411 214782
rect 186313 214570 186379 214573
rect 186313 214568 190164 214570
rect 186313 214512 186318 214568
rect 186374 214512 190164 214568
rect 186313 214510 190164 214512
rect 186313 214507 186379 214510
rect 410057 213618 410123 213621
rect 409830 213616 410123 213618
rect 409830 213560 410062 213616
rect 410118 213560 410123 213616
rect 409830 213558 410123 213560
rect 186313 213482 186379 213485
rect 186313 213480 190164 213482
rect 186313 213424 186318 213480
rect 186374 213424 190164 213480
rect 186313 213422 190164 213424
rect 186313 213419 186379 213422
rect 409830 213044 409890 213558
rect 410057 213555 410123 213558
rect 186313 212258 186379 212261
rect 186313 212256 190164 212258
rect 186313 212200 186318 212256
rect 186374 212200 190164 212256
rect 186313 212198 190164 212200
rect 186313 212195 186379 212198
rect 411437 211170 411503 211173
rect 409860 211168 411503 211170
rect 409860 211112 411442 211168
rect 411498 211112 411503 211168
rect 409860 211110 411503 211112
rect 411437 211107 411503 211110
rect 186405 211034 186471 211037
rect 186405 211032 190164 211034
rect 186405 210976 186410 211032
rect 186466 210976 190164 211032
rect 186405 210974 190164 210976
rect 186405 210971 186471 210974
rect 186313 209946 186379 209949
rect 186313 209944 190164 209946
rect 186313 209888 186318 209944
rect 186374 209888 190164 209944
rect 186313 209886 190164 209888
rect 186313 209883 186379 209886
rect 409873 209538 409939 209541
rect 409830 209536 409939 209538
rect 409830 209480 409878 209536
rect 409934 209480 409939 209536
rect 409830 209475 409939 209480
rect 409830 209236 409890 209475
rect 186957 208722 187023 208725
rect 186957 208720 190164 208722
rect 186957 208664 186962 208720
rect 187018 208664 190164 208720
rect 186957 208662 190164 208664
rect 186957 208659 187023 208662
rect 186313 207634 186379 207637
rect 186313 207632 190164 207634
rect 186313 207576 186318 207632
rect 186374 207576 190164 207632
rect 186313 207574 190164 207576
rect 186313 207571 186379 207574
rect 411253 207362 411319 207365
rect 409860 207360 411319 207362
rect 409860 207304 411258 207360
rect 411314 207304 411319 207360
rect 409860 207302 411319 207304
rect 411253 207299 411319 207302
rect 186313 206410 186379 206413
rect 186313 206408 190164 206410
rect 186313 206352 186318 206408
rect 186374 206352 190164 206408
rect 186313 206350 190164 206352
rect 186313 206347 186379 206350
rect 409321 205594 409387 205597
rect 409321 205592 409522 205594
rect 409321 205536 409326 205592
rect 409382 205536 409522 205592
rect 583520 205580 584960 205820
rect 409321 205534 409522 205536
rect 409321 205531 409387 205534
rect 409462 205428 409522 205534
rect 186313 205322 186379 205325
rect 186313 205320 190164 205322
rect 186313 205264 186318 205320
rect 186374 205264 190164 205320
rect 186313 205262 190164 205264
rect 186313 205259 186379 205262
rect 186405 204098 186471 204101
rect 186405 204096 190164 204098
rect 186405 204040 186410 204096
rect 186466 204040 190164 204096
rect 186405 204038 190164 204040
rect 186405 204035 186471 204038
rect 411253 203554 411319 203557
rect 409860 203552 411319 203554
rect 409860 203496 411258 203552
rect 411314 203496 411319 203552
rect 409860 203494 411319 203496
rect 411253 203491 411319 203494
rect 186313 203010 186379 203013
rect 186313 203008 190164 203010
rect 186313 202952 186318 203008
rect 186374 202952 190164 203008
rect 186313 202950 190164 202952
rect 186313 202947 186379 202950
rect -960 201772 480 202012
rect 186313 201786 186379 201789
rect 186313 201784 190164 201786
rect 186313 201728 186318 201784
rect 186374 201728 190164 201784
rect 186313 201726 190164 201728
rect 186313 201723 186379 201726
rect 411253 201650 411319 201653
rect 409860 201648 411319 201650
rect 409860 201592 411258 201648
rect 411314 201592 411319 201648
rect 409860 201590 411319 201592
rect 411253 201587 411319 201590
rect 186313 200562 186379 200565
rect 186313 200560 190164 200562
rect 186313 200504 186318 200560
rect 186374 200504 190164 200560
rect 186313 200502 190164 200504
rect 186313 200499 186379 200502
rect 411253 199746 411319 199749
rect 409860 199744 411319 199746
rect 409860 199688 411258 199744
rect 411314 199688 411319 199744
rect 409860 199686 411319 199688
rect 411253 199683 411319 199686
rect 186313 199474 186379 199477
rect 186313 199472 190164 199474
rect 186313 199416 186318 199472
rect 186374 199416 190164 199472
rect 186313 199414 190164 199416
rect 186313 199411 186379 199414
rect 186313 198250 186379 198253
rect 186313 198248 190164 198250
rect 186313 198192 186318 198248
rect 186374 198192 190164 198248
rect 186313 198190 190164 198192
rect 186313 198187 186379 198190
rect 411253 197842 411319 197845
rect 409860 197840 411319 197842
rect 409860 197784 411258 197840
rect 411314 197784 411319 197840
rect 409860 197782 411319 197784
rect 411253 197779 411319 197782
rect 187049 197162 187115 197165
rect 187049 197160 190164 197162
rect 187049 197104 187054 197160
rect 187110 197104 190164 197160
rect 187049 197102 190164 197104
rect 187049 197099 187115 197102
rect 186405 195938 186471 195941
rect 411989 195938 412055 195941
rect 186405 195936 190164 195938
rect 186405 195880 186410 195936
rect 186466 195880 190164 195936
rect 186405 195878 190164 195880
rect 409860 195936 412055 195938
rect 409860 195880 411994 195936
rect 412050 195880 412055 195936
rect 409860 195878 412055 195880
rect 186405 195875 186471 195878
rect 411989 195875 412055 195878
rect 186313 194850 186379 194853
rect 186313 194848 190164 194850
rect 186313 194792 186318 194848
rect 186374 194792 190164 194848
rect 186313 194790 190164 194792
rect 186313 194787 186379 194790
rect 411253 194034 411319 194037
rect 409860 194032 411319 194034
rect 409860 193976 411258 194032
rect 411314 193976 411319 194032
rect 409860 193974 411319 193976
rect 411253 193971 411319 193974
rect 186313 193626 186379 193629
rect 186313 193624 190164 193626
rect 186313 193568 186318 193624
rect 186374 193568 190164 193624
rect 186313 193566 190164 193568
rect 186313 193563 186379 193566
rect 186313 192402 186379 192405
rect 186313 192400 190164 192402
rect 186313 192344 186318 192400
rect 186374 192344 190164 192400
rect 583520 192388 584960 192628
rect 186313 192342 190164 192344
rect 186313 192339 186379 192342
rect 411897 192130 411963 192133
rect 409860 192128 411963 192130
rect 409860 192072 411902 192128
rect 411958 192072 411963 192128
rect 409860 192070 411963 192072
rect 411897 192067 411963 192070
rect 186313 191314 186379 191317
rect 186313 191312 190164 191314
rect 186313 191256 186318 191312
rect 186374 191256 190164 191312
rect 186313 191254 190164 191256
rect 186313 191251 186379 191254
rect 411253 190226 411319 190229
rect 409860 190224 411319 190226
rect 409860 190168 411258 190224
rect 411314 190168 411319 190224
rect 409860 190166 411319 190168
rect 411253 190163 411319 190166
rect 186313 190090 186379 190093
rect 186313 190088 190164 190090
rect 186313 190032 186318 190088
rect 186374 190032 190164 190088
rect 186313 190030 190164 190032
rect 186313 190027 186379 190030
rect 186405 189002 186471 189005
rect 186405 189000 190164 189002
rect -960 188716 480 188956
rect 186405 188944 186410 189000
rect 186466 188944 190164 189000
rect 186405 188942 190164 188944
rect 186405 188939 186471 188942
rect 411253 188322 411319 188325
rect 409860 188320 411319 188322
rect 409860 188264 411258 188320
rect 411314 188264 411319 188320
rect 409860 188262 411319 188264
rect 411253 188259 411319 188262
rect 186313 187778 186379 187781
rect 186313 187776 190164 187778
rect 186313 187720 186318 187776
rect 186374 187720 190164 187776
rect 186313 187718 190164 187720
rect 186313 187715 186379 187718
rect 186313 186690 186379 186693
rect 186313 186688 190164 186690
rect 186313 186632 186318 186688
rect 186374 186632 190164 186688
rect 186313 186630 190164 186632
rect 186313 186627 186379 186630
rect 411253 186418 411319 186421
rect 409860 186416 411319 186418
rect 409860 186360 411258 186416
rect 411314 186360 411319 186416
rect 409860 186358 411319 186360
rect 411253 186355 411319 186358
rect 186313 185466 186379 185469
rect 186313 185464 190164 185466
rect 186313 185408 186318 185464
rect 186374 185408 190164 185464
rect 186313 185406 190164 185408
rect 186313 185403 186379 185406
rect 411253 184514 411319 184517
rect 409860 184512 411319 184514
rect 409860 184456 411258 184512
rect 411314 184456 411319 184512
rect 409860 184454 411319 184456
rect 411253 184451 411319 184454
rect 186313 184378 186379 184381
rect 186313 184376 190164 184378
rect 186313 184320 186318 184376
rect 186374 184320 190164 184376
rect 186313 184318 190164 184320
rect 186313 184315 186379 184318
rect 186313 183154 186379 183157
rect 186313 183152 190164 183154
rect 186313 183096 186318 183152
rect 186374 183096 190164 183152
rect 186313 183094 190164 183096
rect 186313 183091 186379 183094
rect 411253 182610 411319 182613
rect 409860 182608 411319 182610
rect 409860 182552 411258 182608
rect 411314 182552 411319 182608
rect 409860 182550 411319 182552
rect 411253 182547 411319 182550
rect 186405 181930 186471 181933
rect 186405 181928 190164 181930
rect 186405 181872 186410 181928
rect 186466 181872 190164 181928
rect 186405 181870 190164 181872
rect 186405 181867 186471 181870
rect 186313 180842 186379 180845
rect 186313 180840 190164 180842
rect 186313 180784 186318 180840
rect 186374 180784 190164 180840
rect 186313 180782 190164 180784
rect 186313 180779 186379 180782
rect 411253 180706 411319 180709
rect 409860 180704 411319 180706
rect 409860 180648 411258 180704
rect 411314 180648 411319 180704
rect 409860 180646 411319 180648
rect 411253 180643 411319 180646
rect 186313 179618 186379 179621
rect 186313 179616 190164 179618
rect 186313 179560 186318 179616
rect 186374 179560 190164 179616
rect 186313 179558 190164 179560
rect 186313 179555 186379 179558
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 411253 178802 411319 178805
rect 409860 178800 411319 178802
rect 409860 178744 411258 178800
rect 411314 178744 411319 178800
rect 409860 178742 411319 178744
rect 411253 178739 411319 178742
rect 186313 178530 186379 178533
rect 186313 178528 190164 178530
rect 186313 178472 186318 178528
rect 186374 178472 190164 178528
rect 186313 178470 190164 178472
rect 186313 178467 186379 178470
rect 186313 177306 186379 177309
rect 186313 177304 190164 177306
rect 186313 177248 186318 177304
rect 186374 177248 190164 177304
rect 186313 177246 190164 177248
rect 186313 177243 186379 177246
rect 411253 177034 411319 177037
rect 409860 177032 411319 177034
rect 409860 176976 411258 177032
rect 411314 176976 411319 177032
rect 409860 176974 411319 176976
rect 411253 176971 411319 176974
rect 186313 176218 186379 176221
rect 186313 176216 190164 176218
rect 186313 176160 186318 176216
rect 186374 176160 190164 176216
rect 186313 176158 190164 176160
rect 186313 176155 186379 176158
rect -960 175796 480 176036
rect 411253 175130 411319 175133
rect 409860 175128 411319 175130
rect 409860 175072 411258 175128
rect 411314 175072 411319 175128
rect 409860 175070 411319 175072
rect 411253 175067 411319 175070
rect 186313 174994 186379 174997
rect 186313 174992 190164 174994
rect 186313 174936 186318 174992
rect 186374 174936 190164 174992
rect 186313 174934 190164 174936
rect 186313 174931 186379 174934
rect 186405 173770 186471 173773
rect 186405 173768 190164 173770
rect 186405 173712 186410 173768
rect 186466 173712 190164 173768
rect 186405 173710 190164 173712
rect 186405 173707 186471 173710
rect 411253 173226 411319 173229
rect 409860 173224 411319 173226
rect 409860 173168 411258 173224
rect 411314 173168 411319 173224
rect 409860 173166 411319 173168
rect 411253 173163 411319 173166
rect 186313 172682 186379 172685
rect 186313 172680 190164 172682
rect 186313 172624 186318 172680
rect 186374 172624 190164 172680
rect 186313 172622 190164 172624
rect 186313 172619 186379 172622
rect 186313 171458 186379 171461
rect 186313 171456 190164 171458
rect 186313 171400 186318 171456
rect 186374 171400 190164 171456
rect 186313 171398 190164 171400
rect 186313 171395 186379 171398
rect 411253 171322 411319 171325
rect 409860 171320 411319 171322
rect 409860 171264 411258 171320
rect 411314 171264 411319 171320
rect 409860 171262 411319 171264
rect 411253 171259 411319 171262
rect 186313 170370 186379 170373
rect 186313 170368 190164 170370
rect 186313 170312 186318 170368
rect 186374 170312 190164 170368
rect 186313 170310 190164 170312
rect 186313 170307 186379 170310
rect 411253 169418 411319 169421
rect 409860 169416 411319 169418
rect 409860 169360 411258 169416
rect 411314 169360 411319 169416
rect 409860 169358 411319 169360
rect 411253 169355 411319 169358
rect 186313 169146 186379 169149
rect 186313 169144 190164 169146
rect 186313 169088 186318 169144
rect 186374 169088 190164 169144
rect 186313 169086 190164 169088
rect 186313 169083 186379 169086
rect 186313 168058 186379 168061
rect 186313 168056 190164 168058
rect 186313 168000 186318 168056
rect 186374 168000 190164 168056
rect 186313 167998 190164 168000
rect 186313 167995 186379 167998
rect 411253 167514 411319 167517
rect 409860 167512 411319 167514
rect 409860 167456 411258 167512
rect 411314 167456 411319 167512
rect 409860 167454 411319 167456
rect 411253 167451 411319 167454
rect 186405 166834 186471 166837
rect 186405 166832 190164 166834
rect 186405 166776 186410 166832
rect 186466 166776 190164 166832
rect 186405 166774 190164 166776
rect 186405 166771 186471 166774
rect 186313 165746 186379 165749
rect 186313 165744 190164 165746
rect 186313 165688 186318 165744
rect 186374 165688 190164 165744
rect 583520 165732 584960 165972
rect 186313 165686 190164 165688
rect 186313 165683 186379 165686
rect 411253 165610 411319 165613
rect 409860 165608 411319 165610
rect 409860 165552 411258 165608
rect 411314 165552 411319 165608
rect 409860 165550 411319 165552
rect 411253 165547 411319 165550
rect 186313 164522 186379 164525
rect 186313 164520 190164 164522
rect 186313 164464 186318 164520
rect 186374 164464 190164 164520
rect 186313 164462 190164 164464
rect 186313 164459 186379 164462
rect 411253 163706 411319 163709
rect 409860 163704 411319 163706
rect 409860 163648 411258 163704
rect 411314 163648 411319 163704
rect 409860 163646 411319 163648
rect 411253 163643 411319 163646
rect 186313 163298 186379 163301
rect 186313 163296 190164 163298
rect 186313 163240 186318 163296
rect 186374 163240 190164 163296
rect 186313 163238 190164 163240
rect 186313 163235 186379 163238
rect -960 162740 480 162980
rect 186313 162210 186379 162213
rect 186313 162208 190164 162210
rect 186313 162152 186318 162208
rect 186374 162152 190164 162208
rect 186313 162150 190164 162152
rect 186313 162147 186379 162150
rect 411253 161802 411319 161805
rect 409860 161800 411319 161802
rect 409860 161744 411258 161800
rect 411314 161744 411319 161800
rect 409860 161742 411319 161744
rect 411253 161739 411319 161742
rect 186313 160986 186379 160989
rect 186313 160984 190164 160986
rect 186313 160928 186318 160984
rect 186374 160928 190164 160984
rect 186313 160926 190164 160928
rect 186313 160923 186379 160926
rect 186313 159898 186379 159901
rect 411253 159898 411319 159901
rect 186313 159896 190164 159898
rect 186313 159840 186318 159896
rect 186374 159840 190164 159896
rect 186313 159838 190164 159840
rect 409860 159896 411319 159898
rect 409860 159840 411258 159896
rect 411314 159840 411319 159896
rect 409860 159838 411319 159840
rect 186313 159835 186379 159838
rect 411253 159835 411319 159838
rect 186405 158674 186471 158677
rect 186405 158672 190164 158674
rect 186405 158616 186410 158672
rect 186466 158616 190164 158672
rect 186405 158614 190164 158616
rect 186405 158611 186471 158614
rect 411253 157994 411319 157997
rect 409860 157992 411319 157994
rect 409860 157936 411258 157992
rect 411314 157936 411319 157992
rect 409860 157934 411319 157936
rect 411253 157931 411319 157934
rect 186313 157586 186379 157589
rect 186313 157584 190164 157586
rect 186313 157528 186318 157584
rect 186374 157528 190164 157584
rect 186313 157526 190164 157528
rect 186313 157523 186379 157526
rect 186313 156362 186379 156365
rect 186313 156360 190164 156362
rect 186313 156304 186318 156360
rect 186374 156304 190164 156360
rect 186313 156302 190164 156304
rect 186313 156299 186379 156302
rect 411253 156090 411319 156093
rect 409860 156088 411319 156090
rect 409860 156032 411258 156088
rect 411314 156032 411319 156088
rect 409860 156030 411319 156032
rect 411253 156027 411319 156030
rect 186313 155274 186379 155277
rect 186313 155272 190164 155274
rect 186313 155216 186318 155272
rect 186374 155216 190164 155272
rect 186313 155214 190164 155216
rect 186313 155211 186379 155214
rect 411253 154186 411319 154189
rect 409860 154184 411319 154186
rect 409860 154128 411258 154184
rect 411314 154128 411319 154184
rect 409860 154126 411319 154128
rect 411253 154123 411319 154126
rect 186313 154050 186379 154053
rect 186313 154048 190164 154050
rect 186313 153992 186318 154048
rect 186374 153992 190164 154048
rect 186313 153990 190164 153992
rect 186313 153987 186379 153990
rect 186313 152826 186379 152829
rect 186313 152824 190164 152826
rect 186313 152768 186318 152824
rect 186374 152768 190164 152824
rect 186313 152766 190164 152768
rect 186313 152763 186379 152766
rect 583520 152540 584960 152780
rect 411253 152282 411319 152285
rect 409860 152280 411319 152282
rect 409860 152224 411258 152280
rect 411314 152224 411319 152280
rect 409860 152222 411319 152224
rect 411253 152219 411319 152222
rect 186405 151738 186471 151741
rect 186405 151736 190164 151738
rect 186405 151680 186410 151736
rect 186466 151680 190164 151736
rect 186405 151678 190164 151680
rect 186405 151675 186471 151678
rect 186313 150514 186379 150517
rect 186313 150512 190164 150514
rect 186313 150456 186318 150512
rect 186374 150456 190164 150512
rect 186313 150454 190164 150456
rect 186313 150451 186379 150454
rect 411253 150378 411319 150381
rect 409860 150376 411319 150378
rect 409860 150320 411258 150376
rect 411314 150320 411319 150376
rect 409860 150318 411319 150320
rect 411253 150315 411319 150318
rect -960 149684 480 149924
rect 186313 149426 186379 149429
rect 186313 149424 190164 149426
rect 186313 149368 186318 149424
rect 186374 149368 190164 149424
rect 186313 149366 190164 149368
rect 186313 149363 186379 149366
rect 411253 148474 411319 148477
rect 409860 148472 411319 148474
rect 409860 148416 411258 148472
rect 411314 148416 411319 148472
rect 409860 148414 411319 148416
rect 411253 148411 411319 148414
rect 186313 148202 186379 148205
rect 186313 148200 190164 148202
rect 186313 148144 186318 148200
rect 186374 148144 190164 148200
rect 186313 148142 190164 148144
rect 186313 148139 186379 148142
rect 186313 147114 186379 147117
rect 186313 147112 190164 147114
rect 186313 147056 186318 147112
rect 186374 147056 190164 147112
rect 186313 147054 190164 147056
rect 186313 147051 186379 147054
rect 411253 146570 411319 146573
rect 409860 146568 411319 146570
rect 409860 146512 411258 146568
rect 411314 146512 411319 146568
rect 409860 146510 411319 146512
rect 411253 146507 411319 146510
rect 186313 145890 186379 145893
rect 186313 145888 190164 145890
rect 186313 145832 186318 145888
rect 186374 145832 190164 145888
rect 186313 145830 190164 145832
rect 186313 145827 186379 145830
rect 186405 144666 186471 144669
rect 411253 144666 411319 144669
rect 186405 144664 190164 144666
rect 186405 144608 186410 144664
rect 186466 144608 190164 144664
rect 186405 144606 190164 144608
rect 409860 144664 411319 144666
rect 409860 144608 411258 144664
rect 411314 144608 411319 144664
rect 409860 144606 411319 144608
rect 186405 144603 186471 144606
rect 411253 144603 411319 144606
rect 186313 143578 186379 143581
rect 186313 143576 190164 143578
rect 186313 143520 186318 143576
rect 186374 143520 190164 143576
rect 186313 143518 190164 143520
rect 186313 143515 186379 143518
rect 411253 142762 411319 142765
rect 409860 142760 411319 142762
rect 409860 142704 411258 142760
rect 411314 142704 411319 142760
rect 409860 142702 411319 142704
rect 411253 142699 411319 142702
rect 186313 142354 186379 142357
rect 186313 142352 190164 142354
rect 186313 142296 186318 142352
rect 186374 142296 190164 142352
rect 186313 142294 190164 142296
rect 186313 142291 186379 142294
rect 187141 141266 187207 141269
rect 187141 141264 190164 141266
rect 187141 141208 187146 141264
rect 187202 141208 190164 141264
rect 187141 141206 190164 141208
rect 187141 141203 187207 141206
rect 411253 140994 411319 140997
rect 409860 140992 411319 140994
rect 409860 140936 411258 140992
rect 411314 140936 411319 140992
rect 409860 140934 411319 140936
rect 411253 140931 411319 140934
rect 186313 140042 186379 140045
rect 186313 140040 190164 140042
rect 186313 139984 186318 140040
rect 186374 139984 190164 140040
rect 186313 139982 190164 139984
rect 186313 139979 186379 139982
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 411253 139090 411319 139093
rect 409860 139088 411319 139090
rect 409860 139032 411258 139088
rect 411314 139032 411319 139088
rect 409860 139030 411319 139032
rect 411253 139027 411319 139030
rect 186313 138954 186379 138957
rect 186313 138952 190164 138954
rect 186313 138896 186318 138952
rect 186374 138896 190164 138952
rect 186313 138894 190164 138896
rect 186313 138891 186379 138894
rect 186313 137730 186379 137733
rect 186313 137728 190164 137730
rect 186313 137672 186318 137728
rect 186374 137672 190164 137728
rect 186313 137670 190164 137672
rect 186313 137667 186379 137670
rect 411253 137186 411319 137189
rect 409860 137184 411319 137186
rect 409860 137128 411258 137184
rect 411314 137128 411319 137184
rect 409860 137126 411319 137128
rect 411253 137123 411319 137126
rect -960 136628 480 136868
rect 186405 136642 186471 136645
rect 186405 136640 190164 136642
rect 186405 136584 186410 136640
rect 186466 136584 190164 136640
rect 186405 136582 190164 136584
rect 186405 136579 186471 136582
rect 186313 135418 186379 135421
rect 186313 135416 190164 135418
rect 186313 135360 186318 135416
rect 186374 135360 190164 135416
rect 186313 135358 190164 135360
rect 186313 135355 186379 135358
rect 411253 135282 411319 135285
rect 409860 135280 411319 135282
rect 409860 135224 411258 135280
rect 411314 135224 411319 135280
rect 409860 135222 411319 135224
rect 411253 135219 411319 135222
rect 187233 134194 187299 134197
rect 187233 134192 190164 134194
rect 187233 134136 187238 134192
rect 187294 134136 190164 134192
rect 187233 134134 190164 134136
rect 187233 134131 187299 134134
rect 411253 133378 411319 133381
rect 409860 133376 411319 133378
rect 409860 133320 411258 133376
rect 411314 133320 411319 133376
rect 409860 133318 411319 133320
rect 411253 133315 411319 133318
rect 186313 133106 186379 133109
rect 186313 133104 190164 133106
rect 186313 133048 186318 133104
rect 186374 133048 190164 133104
rect 186313 133046 190164 133048
rect 186313 133043 186379 133046
rect 186313 131882 186379 131885
rect 186313 131880 190164 131882
rect 186313 131824 186318 131880
rect 186374 131824 190164 131880
rect 186313 131822 190164 131824
rect 186313 131819 186379 131822
rect 411253 131474 411319 131477
rect 409860 131472 411319 131474
rect 409860 131416 411258 131472
rect 411314 131416 411319 131472
rect 409860 131414 411319 131416
rect 411253 131411 411319 131414
rect 186313 130794 186379 130797
rect 186313 130792 190164 130794
rect 186313 130736 186318 130792
rect 186374 130736 190164 130792
rect 186313 130734 190164 130736
rect 186313 130731 186379 130734
rect 129598 129782 130210 129842
rect 129598 129676 129658 129782
rect 130150 129706 130210 129782
rect 131113 129706 131179 129709
rect 130150 129704 131179 129706
rect 130150 129648 131118 129704
rect 131174 129648 131179 129704
rect 130150 129646 131179 129648
rect 131113 129643 131179 129646
rect 186405 129570 186471 129573
rect 411253 129570 411319 129573
rect 186405 129568 190164 129570
rect 186405 129512 186410 129568
rect 186466 129512 190164 129568
rect 186405 129510 190164 129512
rect 409860 129568 411319 129570
rect 409860 129512 411258 129568
rect 411314 129512 411319 129568
rect 409860 129510 411319 129512
rect 186405 129507 186471 129510
rect 411253 129507 411319 129510
rect 131205 129162 131271 129165
rect 130518 129160 131271 129162
rect 130518 129134 131210 129160
rect 129904 129104 131210 129134
rect 131266 129104 131271 129160
rect 129904 129102 131271 129104
rect 129904 129074 130578 129102
rect 131205 129099 131271 129102
rect 437473 128754 437539 128757
rect 440006 128754 440066 129132
rect 437473 128752 440066 128754
rect 437473 128696 437478 128752
rect 437534 128696 440066 128752
rect 437473 128694 440066 128696
rect 437473 128691 437539 128694
rect 131297 128618 131363 128621
rect 130518 128616 131363 128618
rect 130518 128590 131302 128616
rect 129904 128560 131302 128590
rect 131358 128560 131363 128616
rect 129904 128558 131363 128560
rect 129904 128530 130578 128558
rect 131297 128555 131363 128558
rect 186313 128482 186379 128485
rect 186313 128480 190164 128482
rect 186313 128424 186318 128480
rect 186374 128424 190164 128480
rect 186313 128422 190164 128424
rect 186313 128419 186379 128422
rect 132217 127938 132283 127941
rect 130518 127936 132283 127938
rect 130518 127910 132222 127936
rect 129904 127880 132222 127910
rect 132278 127880 132283 127936
rect 129904 127878 132283 127880
rect 129904 127850 130578 127878
rect 132217 127875 132283 127878
rect 411253 127666 411319 127669
rect 409860 127664 411319 127666
rect 409860 127608 411258 127664
rect 411314 127608 411319 127664
rect 409860 127606 411319 127608
rect 411253 127603 411319 127606
rect 132033 127394 132099 127397
rect 130518 127392 132099 127394
rect 130518 127366 132038 127392
rect 129904 127336 132038 127366
rect 132094 127336 132099 127392
rect 129904 127334 132099 127336
rect 129904 127306 130578 127334
rect 132033 127331 132099 127334
rect 186313 127258 186379 127261
rect 186313 127256 190164 127258
rect 186313 127200 186318 127256
rect 186374 127200 190164 127256
rect 186313 127198 190164 127200
rect 186313 127195 186379 127198
rect 437473 127122 437539 127125
rect 440006 127122 440066 127500
rect 437473 127120 440066 127122
rect 437473 127064 437478 127120
rect 437534 127064 440066 127120
rect 437473 127062 440066 127064
rect 437473 127059 437539 127062
rect 131205 126850 131271 126853
rect 130518 126848 131271 126850
rect 130518 126822 131210 126848
rect 129904 126792 131210 126822
rect 131266 126792 131271 126848
rect 129904 126790 131271 126792
rect 129904 126762 130578 126790
rect 131205 126787 131271 126790
rect 131113 126170 131179 126173
rect 130518 126168 131179 126170
rect 130518 126142 131118 126168
rect 129904 126112 131118 126142
rect 131174 126112 131179 126168
rect 129904 126110 131179 126112
rect 129904 126082 130578 126110
rect 131113 126107 131179 126110
rect 186313 126034 186379 126037
rect 539317 126034 539383 126037
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 186313 126032 190164 126034
rect 186313 125976 186318 126032
rect 186374 125976 190164 126032
rect 186313 125974 190164 125976
rect 539317 126032 539426 126034
rect 539317 125976 539322 126032
rect 539378 125976 539426 126032
rect 186313 125971 186379 125974
rect 539317 125971 539426 125976
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 411253 125762 411319 125765
rect 409860 125760 411319 125762
rect 409860 125704 411258 125760
rect 411314 125704 411319 125760
rect 409860 125702 411319 125704
rect 411253 125699 411319 125702
rect 437473 125762 437539 125765
rect 440006 125762 440066 125868
rect 437473 125760 440066 125762
rect 437473 125704 437478 125760
rect 437534 125704 440066 125760
rect 437473 125702 440066 125704
rect 437473 125699 437539 125702
rect 132033 125626 132099 125629
rect 130150 125624 132099 125626
rect 130150 125592 132038 125624
rect 129904 125568 132038 125592
rect 132094 125568 132099 125624
rect 129904 125566 132099 125568
rect 129904 125532 130210 125566
rect 132033 125563 132099 125566
rect 539366 125460 539426 125971
rect 583520 125884 584960 125974
rect 131113 125082 131179 125085
rect 130518 125080 131179 125082
rect 130518 125054 131118 125080
rect 129904 125024 131118 125054
rect 131174 125024 131179 125080
rect 129904 125022 131179 125024
rect 129904 124994 130578 125022
rect 131113 125019 131179 125022
rect 186313 124946 186379 124949
rect 186313 124944 190164 124946
rect 186313 124888 186318 124944
rect 186374 124888 190164 124944
rect 186313 124886 190164 124888
rect 186313 124883 186379 124886
rect 131205 124538 131271 124541
rect 130518 124536 131271 124538
rect 130518 124510 131210 124536
rect 129904 124480 131210 124510
rect 131266 124480 131271 124536
rect 129904 124478 131271 124480
rect 129904 124450 130578 124478
rect 131205 124475 131271 124478
rect 437473 124402 437539 124405
rect 437473 124400 440066 124402
rect 437473 124344 437478 124400
rect 437534 124344 440066 124400
rect 437473 124342 440066 124344
rect 437473 124339 437539 124342
rect 440006 124236 440066 124342
rect 132217 123858 132283 123861
rect 411253 123858 411319 123861
rect 130518 123856 132283 123858
rect 130518 123830 132222 123856
rect -960 123572 480 123812
rect 129904 123800 132222 123830
rect 132278 123800 132283 123856
rect 129904 123798 132283 123800
rect 409860 123856 411319 123858
rect 409860 123800 411258 123856
rect 411314 123800 411319 123856
rect 409860 123798 411319 123800
rect 129904 123770 130578 123798
rect 132217 123795 132283 123798
rect 411253 123795 411319 123798
rect 187325 123722 187391 123725
rect 187325 123720 190164 123722
rect 187325 123664 187330 123720
rect 187386 123664 190164 123720
rect 187325 123662 190164 123664
rect 187325 123659 187391 123662
rect 131113 123314 131179 123317
rect 130518 123312 131179 123314
rect 130518 123286 131118 123312
rect 129904 123256 131118 123286
rect 131174 123256 131179 123312
rect 129904 123254 131179 123256
rect 129904 123226 130578 123254
rect 131113 123251 131179 123254
rect 131205 122770 131271 122773
rect 130518 122768 131271 122770
rect 130518 122742 131210 122768
rect 129904 122712 131210 122742
rect 131266 122712 131271 122768
rect 129904 122710 131271 122712
rect 129904 122682 130578 122710
rect 131205 122707 131271 122710
rect 186313 122634 186379 122637
rect 186313 122632 190164 122634
rect 186313 122576 186318 122632
rect 186374 122576 190164 122632
rect 186313 122574 190164 122576
rect 186313 122571 186379 122574
rect 131205 122090 131271 122093
rect 130518 122088 131271 122090
rect 130518 122062 131210 122088
rect 129904 122032 131210 122062
rect 131266 122032 131271 122088
rect 129904 122030 131271 122032
rect 129904 122002 130578 122030
rect 131205 122027 131271 122030
rect 411253 121954 411319 121957
rect 409860 121952 411319 121954
rect 409860 121896 411258 121952
rect 411314 121896 411319 121952
rect 409860 121894 411319 121896
rect 411253 121891 411319 121894
rect 437473 121954 437539 121957
rect 440006 121954 440066 122468
rect 437473 121952 440066 121954
rect 437473 121896 437478 121952
rect 437534 121896 440066 121952
rect 437473 121894 440066 121896
rect 437473 121891 437539 121894
rect 131113 121546 131179 121549
rect 130518 121544 131179 121546
rect 130518 121518 131118 121544
rect 129904 121488 131118 121518
rect 131174 121488 131179 121544
rect 129904 121486 131179 121488
rect 129904 121458 130578 121486
rect 131113 121483 131179 121486
rect 186405 121410 186471 121413
rect 186405 121408 190164 121410
rect 186405 121352 186410 121408
rect 186466 121352 190164 121408
rect 186405 121350 190164 121352
rect 186405 121347 186471 121350
rect 131205 121002 131271 121005
rect 130518 121000 131271 121002
rect 130518 120974 131210 121000
rect 129904 120944 131210 120974
rect 131266 120944 131271 121000
rect 129904 120942 131271 120944
rect 129904 120914 130578 120942
rect 131205 120939 131271 120942
rect 437473 120458 437539 120461
rect 440006 120458 440066 120836
rect 437473 120456 440066 120458
rect 437473 120400 437478 120456
rect 437534 120400 440066 120456
rect 437473 120398 440066 120400
rect 437473 120395 437539 120398
rect 131941 120322 132007 120325
rect 130518 120320 132007 120322
rect 130518 120294 131946 120320
rect 129904 120264 131946 120294
rect 132002 120264 132007 120320
rect 129904 120262 132007 120264
rect 129904 120234 130578 120262
rect 131941 120259 132007 120262
rect 186313 120322 186379 120325
rect 186313 120320 190164 120322
rect 186313 120264 186318 120320
rect 186374 120264 190164 120320
rect 186313 120262 190164 120264
rect 186313 120259 186379 120262
rect 411253 120050 411319 120053
rect 409860 120048 411319 120050
rect 409860 119992 411258 120048
rect 411314 119992 411319 120048
rect 409860 119990 411319 119992
rect 411253 119987 411319 119990
rect 132217 119778 132283 119781
rect 130518 119776 132283 119778
rect 130518 119750 132222 119776
rect 129904 119720 132222 119750
rect 132278 119720 132283 119776
rect 129904 119718 132283 119720
rect 129904 119690 130578 119718
rect 132217 119715 132283 119718
rect 437565 119642 437631 119645
rect 437565 119640 440066 119642
rect 437565 119584 437570 119640
rect 437626 119584 440066 119640
rect 437565 119582 440066 119584
rect 437565 119579 437631 119582
rect 131113 119234 131179 119237
rect 130518 119232 131179 119234
rect 130518 119206 131118 119232
rect 129904 119176 131118 119206
rect 131174 119176 131179 119232
rect 440006 119204 440066 119582
rect 129904 119174 131179 119176
rect 129904 119146 130578 119174
rect 131113 119171 131179 119174
rect 186313 119098 186379 119101
rect 186313 119096 190164 119098
rect 186313 119040 186318 119096
rect 186374 119040 190164 119096
rect 186313 119038 190164 119040
rect 186313 119035 186379 119038
rect 131205 118690 131271 118693
rect 130518 118688 131271 118690
rect 130518 118662 131210 118688
rect 129904 118632 131210 118662
rect 131266 118632 131271 118688
rect 129904 118630 131271 118632
rect 129904 118602 130578 118630
rect 131205 118627 131271 118630
rect 411253 118146 411319 118149
rect 409860 118144 411319 118146
rect 409860 118088 411258 118144
rect 411314 118088 411319 118144
rect 409860 118086 411319 118088
rect 411253 118083 411319 118086
rect 437473 118146 437539 118149
rect 437473 118144 440066 118146
rect 437473 118088 437478 118144
rect 437534 118088 440066 118144
rect 437473 118086 440066 118088
rect 437473 118083 437539 118086
rect 131113 118010 131179 118013
rect 130518 118008 131179 118010
rect 130518 117982 131118 118008
rect 129904 117952 131118 117982
rect 131174 117952 131179 118008
rect 129904 117950 131179 117952
rect 129904 117922 130578 117950
rect 131113 117947 131179 117950
rect 186313 118010 186379 118013
rect 186313 118008 190164 118010
rect 186313 117952 186318 118008
rect 186374 117952 190164 118008
rect 186313 117950 190164 117952
rect 186313 117947 186379 117950
rect 440006 117572 440066 118086
rect 131205 117466 131271 117469
rect 130518 117464 131271 117466
rect 130518 117438 131210 117464
rect 129904 117408 131210 117438
rect 131266 117408 131271 117464
rect 129904 117406 131271 117408
rect 129904 117378 130578 117406
rect 131205 117403 131271 117406
rect 131205 116922 131271 116925
rect 130518 116920 131271 116922
rect 130518 116894 131210 116920
rect 129904 116864 131210 116894
rect 131266 116864 131271 116920
rect 129904 116862 131271 116864
rect 129904 116834 130578 116862
rect 131205 116859 131271 116862
rect 186313 116786 186379 116789
rect 186313 116784 190164 116786
rect 186313 116728 186318 116784
rect 186374 116728 190164 116784
rect 186313 116726 190164 116728
rect 186313 116723 186379 116726
rect 542537 116378 542603 116381
rect 539948 116376 542603 116378
rect 539948 116320 542542 116376
rect 542598 116320 542603 116376
rect 539948 116318 542603 116320
rect 542537 116315 542603 116318
rect 131113 116242 131179 116245
rect 411253 116242 411319 116245
rect 130518 116240 131179 116242
rect 130518 116214 131118 116240
rect 129904 116184 131118 116214
rect 131174 116184 131179 116240
rect 129904 116182 131179 116184
rect 409860 116240 411319 116242
rect 409860 116184 411258 116240
rect 411314 116184 411319 116240
rect 409860 116182 411319 116184
rect 129904 116154 130578 116182
rect 131113 116179 131179 116182
rect 411253 116179 411319 116182
rect 131205 115698 131271 115701
rect 130518 115696 131271 115698
rect 130518 115670 131210 115696
rect 129904 115640 131210 115670
rect 131266 115640 131271 115696
rect 129904 115638 131271 115640
rect 129904 115610 130578 115638
rect 131205 115635 131271 115638
rect 437473 115698 437539 115701
rect 440006 115698 440066 115804
rect 437473 115696 440066 115698
rect 437473 115640 437478 115696
rect 437534 115640 440066 115696
rect 437473 115638 440066 115640
rect 437473 115635 437539 115638
rect 186313 115562 186379 115565
rect 186313 115560 190164 115562
rect 186313 115504 186318 115560
rect 186374 115504 190164 115560
rect 186313 115502 190164 115504
rect 186313 115499 186379 115502
rect 131205 115154 131271 115157
rect 130518 115152 131271 115154
rect 130518 115126 131210 115152
rect 129904 115096 131210 115126
rect 131266 115096 131271 115152
rect 129904 115094 131271 115096
rect 129904 115066 130578 115094
rect 131205 115091 131271 115094
rect 131205 114474 131271 114477
rect 130518 114472 131271 114474
rect 130518 114446 131210 114472
rect 129904 114416 131210 114446
rect 131266 114416 131271 114472
rect 129904 114414 131271 114416
rect 129904 114386 130578 114414
rect 131205 114411 131271 114414
rect 187417 114474 187483 114477
rect 437473 114474 437539 114477
rect 187417 114472 190164 114474
rect 187417 114416 187422 114472
rect 187478 114416 190164 114472
rect 187417 114414 190164 114416
rect 437473 114472 440066 114474
rect 437473 114416 437478 114472
rect 437534 114416 440066 114472
rect 437473 114414 440066 114416
rect 187417 114411 187483 114414
rect 437473 114411 437539 114414
rect 411989 114338 412055 114341
rect 409860 114336 412055 114338
rect 409860 114280 411994 114336
rect 412050 114280 412055 114336
rect 409860 114278 412055 114280
rect 411989 114275 412055 114278
rect 440006 114172 440066 114414
rect 131297 113930 131363 113933
rect 130518 113928 131363 113930
rect 130518 113902 131302 113928
rect 129904 113872 131302 113902
rect 131358 113872 131363 113928
rect 129904 113870 131363 113872
rect 129904 113842 130578 113870
rect 131297 113867 131363 113870
rect 131113 113386 131179 113389
rect 130518 113384 131179 113386
rect 130518 113358 131118 113384
rect 129904 113328 131118 113358
rect 131174 113328 131179 113384
rect 129904 113326 131179 113328
rect 129904 113298 130578 113326
rect 131113 113323 131179 113326
rect 186957 113250 187023 113253
rect 186957 113248 190164 113250
rect 186957 113192 186962 113248
rect 187018 113192 190164 113248
rect 186957 113190 190164 113192
rect 186957 113187 187023 113190
rect 131205 112842 131271 112845
rect 130518 112840 131271 112842
rect 130518 112814 131210 112840
rect 129904 112784 131210 112814
rect 131266 112784 131271 112840
rect 129904 112782 131271 112784
rect 129904 112754 130578 112782
rect 131205 112779 131271 112782
rect 437473 112842 437539 112845
rect 437473 112840 440066 112842
rect 437473 112784 437478 112840
rect 437534 112784 440066 112840
rect 437473 112782 440066 112784
rect 437473 112779 437539 112782
rect 440006 112540 440066 112782
rect 583520 112692 584960 112932
rect 411253 112434 411319 112437
rect 409860 112432 411319 112434
rect 409860 112376 411258 112432
rect 411314 112376 411319 112432
rect 409860 112374 411319 112376
rect 411253 112371 411319 112374
rect 131113 112162 131179 112165
rect 130518 112160 131179 112162
rect 130518 112134 131118 112160
rect 129904 112104 131118 112134
rect 131174 112104 131179 112160
rect 129904 112102 131179 112104
rect 129904 112074 130578 112102
rect 131113 112099 131179 112102
rect 186313 112162 186379 112165
rect 186313 112160 190164 112162
rect 186313 112104 186318 112160
rect 186374 112104 190164 112160
rect 186313 112102 190164 112104
rect 186313 112099 186379 112102
rect 132125 111618 132191 111621
rect 130518 111616 132191 111618
rect 130518 111590 132130 111616
rect 129904 111560 132130 111590
rect 132186 111560 132191 111616
rect 129904 111558 132191 111560
rect 129904 111530 130578 111558
rect 132125 111555 132191 111558
rect 437473 111346 437539 111349
rect 437473 111344 440066 111346
rect 437473 111288 437478 111344
rect 437534 111288 440066 111344
rect 437473 111286 440066 111288
rect 437473 111283 437539 111286
rect 131205 111074 131271 111077
rect 130518 111072 131271 111074
rect 130518 111046 131210 111072
rect 129904 111016 131210 111046
rect 131266 111016 131271 111072
rect 129904 111014 131271 111016
rect 129904 110986 130578 111014
rect 131205 111011 131271 111014
rect 186313 110938 186379 110941
rect 186313 110936 190164 110938
rect 186313 110880 186318 110936
rect 186374 110880 190164 110936
rect 440006 110908 440066 111286
rect 186313 110878 190164 110880
rect 186313 110875 186379 110878
rect -960 110516 480 110756
rect 411253 110530 411319 110533
rect 409860 110528 411319 110530
rect 409860 110472 411258 110528
rect 411314 110472 411319 110528
rect 409860 110470 411319 110472
rect 411253 110467 411319 110470
rect 131205 110394 131271 110397
rect 130518 110392 131271 110394
rect 130518 110366 131210 110392
rect 129904 110336 131210 110366
rect 131266 110336 131271 110392
rect 129904 110334 131271 110336
rect 129904 110306 130578 110334
rect 131205 110331 131271 110334
rect 131113 109850 131179 109853
rect 130518 109848 131179 109850
rect 130518 109822 131118 109848
rect 129904 109792 131118 109822
rect 131174 109792 131179 109848
rect 129904 109790 131179 109792
rect 129904 109762 130578 109790
rect 131113 109787 131179 109790
rect 186313 109850 186379 109853
rect 186313 109848 190164 109850
rect 186313 109792 186318 109848
rect 186374 109792 190164 109848
rect 186313 109790 190164 109792
rect 186313 109787 186379 109790
rect 437473 109714 437539 109717
rect 437473 109712 440066 109714
rect 437473 109656 437478 109712
rect 437534 109656 440066 109712
rect 437473 109654 440066 109656
rect 437473 109651 437539 109654
rect 131297 109306 131363 109309
rect 130518 109304 131363 109306
rect 130518 109278 131302 109304
rect 129904 109248 131302 109278
rect 131358 109248 131363 109304
rect 129904 109246 131363 109248
rect 129904 109218 130578 109246
rect 131297 109243 131363 109246
rect 440006 109140 440066 109654
rect 131205 108626 131271 108629
rect 130518 108624 131271 108626
rect 130518 108598 131210 108624
rect 129904 108568 131210 108598
rect 131266 108568 131271 108624
rect 129904 108566 131271 108568
rect 129904 108538 130578 108566
rect 131205 108563 131271 108566
rect 186313 108626 186379 108629
rect 411897 108626 411963 108629
rect 186313 108624 190164 108626
rect 186313 108568 186318 108624
rect 186374 108568 190164 108624
rect 186313 108566 190164 108568
rect 409860 108624 411963 108626
rect 409860 108568 411902 108624
rect 411958 108568 411963 108624
rect 409860 108566 411963 108568
rect 186313 108563 186379 108566
rect 411897 108563 411963 108566
rect 131113 108082 131179 108085
rect 130518 108080 131179 108082
rect 130518 108054 131118 108080
rect 129904 108024 131118 108054
rect 131174 108024 131179 108080
rect 129904 108022 131179 108024
rect 129904 107994 130578 108022
rect 131113 108019 131179 108022
rect 131205 107538 131271 107541
rect 130518 107536 131271 107538
rect 130518 107510 131210 107536
rect 129904 107480 131210 107510
rect 131266 107480 131271 107536
rect 129904 107478 131271 107480
rect 129904 107450 130578 107478
rect 131205 107475 131271 107478
rect 186405 107538 186471 107541
rect 186405 107536 190164 107538
rect 186405 107480 186410 107536
rect 186466 107480 190164 107536
rect 186405 107478 190164 107480
rect 186405 107475 186471 107478
rect 436737 107402 436803 107405
rect 440006 107402 440066 107508
rect 436737 107400 440066 107402
rect 436737 107344 436742 107400
rect 436798 107344 440066 107400
rect 436737 107342 440066 107344
rect 436737 107339 436803 107342
rect 542445 107266 542511 107269
rect 539948 107264 542511 107266
rect 539948 107208 542450 107264
rect 542506 107208 542511 107264
rect 539948 107206 542511 107208
rect 542445 107203 542511 107206
rect 131113 106994 131179 106997
rect 130518 106992 131179 106994
rect 130518 106966 131118 106992
rect 129904 106936 131118 106966
rect 131174 106936 131179 106992
rect 129904 106934 131179 106936
rect 129904 106906 130578 106934
rect 131113 106931 131179 106934
rect 411253 106722 411319 106725
rect 409860 106720 411319 106722
rect 409860 106664 411258 106720
rect 411314 106664 411319 106720
rect 409860 106662 411319 106664
rect 411253 106659 411319 106662
rect 131297 106314 131363 106317
rect 130150 106312 131363 106314
rect 130150 106280 131302 106312
rect 129904 106256 131302 106280
rect 131358 106256 131363 106312
rect 129904 106254 131363 106256
rect 129904 106220 130210 106254
rect 131297 106251 131363 106254
rect 186313 106314 186379 106317
rect 186313 106312 190164 106314
rect 186313 106256 186318 106312
rect 186374 106256 190164 106312
rect 186313 106254 190164 106256
rect 186313 106251 186379 106254
rect 437473 106042 437539 106045
rect 437473 106040 440066 106042
rect 437473 105984 437478 106040
rect 437534 105984 440066 106040
rect 437473 105982 440066 105984
rect 437473 105979 437539 105982
rect 440006 105876 440066 105982
rect 131113 105770 131179 105773
rect 130518 105768 131179 105770
rect 130518 105742 131118 105768
rect 129904 105712 131118 105742
rect 131174 105712 131179 105768
rect 129904 105710 131179 105712
rect 129904 105682 130578 105710
rect 131113 105707 131179 105710
rect 131205 105226 131271 105229
rect 130518 105224 131271 105226
rect 130518 105198 131210 105224
rect 129904 105168 131210 105198
rect 131266 105168 131271 105224
rect 129904 105166 131271 105168
rect 129904 105138 130578 105166
rect 131205 105163 131271 105166
rect 186313 105090 186379 105093
rect 186313 105088 190164 105090
rect 186313 105032 186318 105088
rect 186374 105032 190164 105088
rect 186313 105030 190164 105032
rect 186313 105027 186379 105030
rect 411253 104818 411319 104821
rect 409860 104816 411319 104818
rect 409860 104760 411258 104816
rect 411314 104760 411319 104816
rect 409860 104758 411319 104760
rect 411253 104755 411319 104758
rect 437657 104818 437723 104821
rect 437657 104816 440066 104818
rect 437657 104760 437662 104816
rect 437718 104760 440066 104816
rect 437657 104758 440066 104760
rect 437657 104755 437723 104758
rect 131205 104546 131271 104549
rect 130518 104544 131271 104546
rect 130518 104518 131210 104544
rect 129904 104488 131210 104518
rect 131266 104488 131271 104544
rect 129904 104486 131271 104488
rect 129904 104458 130578 104486
rect 131205 104483 131271 104486
rect 440006 104244 440066 104758
rect 131113 104002 131179 104005
rect 130518 104000 131179 104002
rect 130518 103974 131118 104000
rect 129904 103944 131118 103974
rect 131174 103944 131179 104000
rect 129904 103942 131179 103944
rect 129904 103914 130578 103942
rect 131113 103939 131179 103942
rect 186313 104002 186379 104005
rect 186313 104000 190164 104002
rect 186313 103944 186318 104000
rect 186374 103944 190164 104000
rect 186313 103942 190164 103944
rect 186313 103939 186379 103942
rect 131205 103458 131271 103461
rect 130518 103456 131271 103458
rect 130518 103430 131210 103456
rect 129904 103400 131210 103430
rect 131266 103400 131271 103456
rect 129904 103398 131271 103400
rect 129904 103370 130578 103398
rect 131205 103395 131271 103398
rect 411253 103050 411319 103053
rect 409860 103048 411319 103050
rect 409860 102992 411258 103048
rect 411314 102992 411319 103048
rect 409860 102990 411319 102992
rect 411253 102987 411319 102990
rect 437473 103050 437539 103053
rect 437473 103048 440066 103050
rect 437473 102992 437478 103048
rect 437534 102992 440066 103048
rect 437473 102990 440066 102992
rect 437473 102987 437539 102990
rect 131665 102778 131731 102781
rect 130518 102776 131731 102778
rect 130518 102750 131670 102776
rect 129904 102720 131670 102750
rect 131726 102720 131731 102776
rect 129904 102718 131731 102720
rect 129904 102690 130578 102718
rect 131665 102715 131731 102718
rect 186313 102778 186379 102781
rect 186313 102776 190164 102778
rect 186313 102720 186318 102776
rect 186374 102720 190164 102776
rect 186313 102718 190164 102720
rect 186313 102715 186379 102718
rect 440006 102476 440066 102990
rect 131113 102234 131179 102237
rect 130518 102232 131179 102234
rect 130518 102206 131118 102232
rect 129904 102176 131118 102206
rect 131174 102176 131179 102232
rect 129904 102174 131179 102176
rect 129904 102146 130578 102174
rect 131113 102171 131179 102174
rect 131205 101690 131271 101693
rect 130518 101688 131271 101690
rect 130518 101662 131210 101688
rect 129904 101632 131210 101662
rect 131266 101632 131271 101688
rect 129904 101630 131271 101632
rect 129904 101602 130578 101630
rect 131205 101627 131271 101630
rect 186313 101690 186379 101693
rect 186313 101688 190164 101690
rect 186313 101632 186318 101688
rect 186374 101632 190164 101688
rect 186313 101630 190164 101632
rect 186313 101627 186379 101630
rect 437473 101418 437539 101421
rect 437473 101416 440066 101418
rect 437473 101360 437478 101416
rect 437534 101360 440066 101416
rect 437473 101358 440066 101360
rect 437473 101355 437539 101358
rect 131113 101146 131179 101149
rect 411253 101146 411319 101149
rect 130518 101144 131179 101146
rect 130518 101118 131118 101144
rect 129904 101088 131118 101118
rect 131174 101088 131179 101144
rect 129904 101086 131179 101088
rect 409860 101144 411319 101146
rect 409860 101088 411258 101144
rect 411314 101088 411319 101144
rect 409860 101086 411319 101088
rect 129904 101058 130578 101086
rect 131113 101083 131179 101086
rect 411253 101083 411319 101086
rect 440006 100844 440066 101358
rect 131849 100466 131915 100469
rect 130518 100464 131915 100466
rect 130518 100438 131854 100464
rect 129904 100408 131854 100438
rect 131910 100408 131915 100464
rect 129904 100406 131915 100408
rect 129904 100378 130578 100406
rect 131849 100403 131915 100406
rect 186313 100466 186379 100469
rect 186313 100464 190164 100466
rect 186313 100408 186318 100464
rect 186374 100408 190164 100464
rect 186313 100406 190164 100408
rect 186313 100403 186379 100406
rect 131205 99922 131271 99925
rect 130518 99920 131271 99922
rect 130518 99894 131210 99920
rect 129904 99864 131210 99894
rect 131266 99864 131271 99920
rect 129904 99862 131271 99864
rect 129904 99834 130578 99862
rect 131205 99859 131271 99862
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 131205 99378 131271 99381
rect 130518 99376 131271 99378
rect 130518 99350 131210 99376
rect 129904 99320 131210 99350
rect 131266 99320 131271 99376
rect 129904 99318 131271 99320
rect 129904 99290 130578 99318
rect 131205 99315 131271 99318
rect 186405 99378 186471 99381
rect 437473 99378 437539 99381
rect 186405 99376 190164 99378
rect 186405 99320 186410 99376
rect 186466 99320 190164 99376
rect 186405 99318 190164 99320
rect 437473 99376 440066 99378
rect 437473 99320 437478 99376
rect 437534 99320 440066 99376
rect 583520 99364 584960 99454
rect 437473 99318 440066 99320
rect 186405 99315 186471 99318
rect 437473 99315 437539 99318
rect 411253 99242 411319 99245
rect 409860 99240 411319 99242
rect 409860 99184 411258 99240
rect 411314 99184 411319 99240
rect 440006 99212 440066 99318
rect 409860 99182 411319 99184
rect 411253 99179 411319 99182
rect 131113 98698 131179 98701
rect 130518 98696 131179 98698
rect 130518 98670 131118 98696
rect 129904 98640 131118 98670
rect 131174 98640 131179 98696
rect 129904 98638 131179 98640
rect 129904 98610 130578 98638
rect 131113 98635 131179 98638
rect 131481 98154 131547 98157
rect 130518 98152 131547 98154
rect 130518 98126 131486 98152
rect 129904 98096 131486 98126
rect 131542 98096 131547 98152
rect 129904 98094 131547 98096
rect 129904 98066 130578 98094
rect 131481 98091 131547 98094
rect 186313 98154 186379 98157
rect 542353 98154 542419 98157
rect 186313 98152 190164 98154
rect 186313 98096 186318 98152
rect 186374 98096 190164 98152
rect 186313 98094 190164 98096
rect 539948 98152 542419 98154
rect 539948 98096 542358 98152
rect 542414 98096 542419 98152
rect 539948 98094 542419 98096
rect 186313 98091 186379 98094
rect 542353 98091 542419 98094
rect 437473 97746 437539 97749
rect 437473 97744 440066 97746
rect -960 97460 480 97700
rect 437473 97688 437478 97744
rect 437534 97688 440066 97744
rect 437473 97686 440066 97688
rect 437473 97683 437539 97686
rect 131205 97610 131271 97613
rect 130518 97608 131271 97610
rect 130518 97582 131210 97608
rect 129904 97552 131210 97582
rect 131266 97552 131271 97608
rect 440006 97580 440066 97686
rect 129904 97550 131271 97552
rect 129904 97522 130578 97550
rect 131205 97547 131271 97550
rect 412081 97338 412147 97341
rect 409860 97336 412147 97338
rect 409860 97280 412086 97336
rect 412142 97280 412147 97336
rect 409860 97278 412147 97280
rect 412081 97275 412147 97278
rect 131113 97066 131179 97069
rect 130518 97064 131179 97066
rect 130518 97038 131118 97064
rect 129904 97008 131118 97038
rect 131174 97008 131179 97064
rect 129904 97006 131179 97008
rect 129904 96978 130578 97006
rect 131113 97003 131179 97006
rect 186313 96930 186379 96933
rect 186313 96928 190164 96930
rect 186313 96872 186318 96928
rect 186374 96872 190164 96928
rect 186313 96870 190164 96872
rect 186313 96867 186379 96870
rect 131205 96386 131271 96389
rect 130518 96384 131271 96386
rect 130518 96358 131210 96384
rect 129904 96328 131210 96358
rect 131266 96328 131271 96384
rect 129904 96326 131271 96328
rect 129904 96298 130578 96326
rect 131205 96323 131271 96326
rect 437473 96250 437539 96253
rect 437473 96248 440066 96250
rect 437473 96192 437478 96248
rect 437534 96192 440066 96248
rect 437473 96190 440066 96192
rect 437473 96187 437539 96190
rect 131113 95842 131179 95845
rect 130518 95840 131179 95842
rect 130518 95814 131118 95840
rect 129904 95784 131118 95814
rect 131174 95784 131179 95840
rect 129904 95782 131179 95784
rect 129904 95754 130578 95782
rect 131113 95779 131179 95782
rect 186313 95842 186379 95845
rect 186313 95840 190164 95842
rect 186313 95784 186318 95840
rect 186374 95784 190164 95840
rect 440006 95812 440066 96190
rect 186313 95782 190164 95784
rect 186313 95779 186379 95782
rect 411805 95434 411871 95437
rect 409860 95432 411871 95434
rect 409860 95376 411810 95432
rect 411866 95376 411871 95432
rect 409860 95374 411871 95376
rect 411805 95371 411871 95374
rect 132217 95298 132283 95301
rect 130518 95296 132283 95298
rect 130518 95270 132222 95296
rect 129904 95240 132222 95270
rect 132278 95240 132283 95296
rect 129904 95238 132283 95240
rect 129904 95210 130578 95238
rect 132217 95235 132283 95238
rect 437473 94754 437539 94757
rect 437473 94752 440066 94754
rect 437473 94696 437478 94752
rect 437534 94696 440066 94752
rect 437473 94694 440066 94696
rect 437473 94691 437539 94694
rect 131205 94618 131271 94621
rect 130518 94616 131271 94618
rect 130518 94590 131210 94616
rect 129904 94560 131210 94590
rect 131266 94560 131271 94616
rect 129904 94558 131271 94560
rect 129904 94530 130578 94558
rect 131205 94555 131271 94558
rect 186313 94618 186379 94621
rect 186313 94616 190164 94618
rect 186313 94560 186318 94616
rect 186374 94560 190164 94616
rect 186313 94558 190164 94560
rect 186313 94555 186379 94558
rect 440006 94180 440066 94694
rect 131113 94074 131179 94077
rect 130518 94072 131179 94074
rect 130518 94046 131118 94072
rect 129904 94016 131118 94046
rect 131174 94016 131179 94072
rect 129904 94014 131179 94016
rect 129904 93986 130578 94014
rect 131113 94011 131179 94014
rect 131205 93530 131271 93533
rect 130518 93528 131271 93530
rect 130518 93502 131210 93528
rect 129904 93472 131210 93502
rect 131266 93472 131271 93528
rect 129904 93470 131271 93472
rect 129904 93442 130578 93470
rect 131205 93467 131271 93470
rect 186313 93530 186379 93533
rect 411345 93530 411411 93533
rect 186313 93528 190164 93530
rect 186313 93472 186318 93528
rect 186374 93472 190164 93528
rect 186313 93470 190164 93472
rect 409860 93528 411411 93530
rect 409860 93472 411350 93528
rect 411406 93472 411411 93528
rect 409860 93470 411411 93472
rect 186313 93467 186379 93470
rect 411345 93467 411411 93470
rect 437473 93122 437539 93125
rect 437473 93120 440066 93122
rect 437473 93064 437478 93120
rect 437534 93064 440066 93120
rect 437473 93062 440066 93064
rect 437473 93059 437539 93062
rect 131113 92850 131179 92853
rect 130518 92848 131179 92850
rect 130518 92822 131118 92848
rect 129904 92792 131118 92822
rect 131174 92792 131179 92848
rect 129904 92790 131179 92792
rect 129904 92762 130578 92790
rect 131113 92787 131179 92790
rect 440006 92548 440066 93062
rect 131205 92306 131271 92309
rect 130518 92304 131271 92306
rect 130518 92278 131210 92304
rect 129904 92248 131210 92278
rect 131266 92248 131271 92304
rect 129904 92246 131271 92248
rect 129904 92218 130578 92246
rect 131205 92243 131271 92246
rect 187509 92306 187575 92309
rect 187509 92304 190164 92306
rect 187509 92248 187514 92304
rect 187570 92248 190164 92304
rect 187509 92246 190164 92248
rect 187509 92243 187575 92246
rect 131113 91762 131179 91765
rect 130518 91760 131179 91762
rect 130518 91734 131118 91760
rect 129904 91704 131118 91734
rect 131174 91704 131179 91760
rect 129904 91702 131179 91704
rect 129904 91674 130578 91702
rect 131113 91699 131179 91702
rect 411253 91626 411319 91629
rect 409860 91624 411319 91626
rect 409860 91568 411258 91624
rect 411314 91568 411319 91624
rect 409860 91566 411319 91568
rect 411253 91563 411319 91566
rect 131297 91218 131363 91221
rect 130518 91216 131363 91218
rect 130518 91190 131302 91216
rect 129904 91160 131302 91190
rect 131358 91160 131363 91216
rect 129904 91158 131363 91160
rect 129904 91130 130578 91158
rect 131297 91155 131363 91158
rect 186313 91218 186379 91221
rect 186313 91216 190164 91218
rect 186313 91160 186318 91216
rect 186374 91160 190164 91216
rect 186313 91158 190164 91160
rect 186313 91155 186379 91158
rect 437473 91082 437539 91085
rect 437473 91080 440066 91082
rect 437473 91024 437478 91080
rect 437534 91024 440066 91080
rect 437473 91022 440066 91024
rect 437473 91019 437539 91022
rect 440006 90916 440066 91022
rect 131205 90538 131271 90541
rect 130518 90536 131271 90538
rect 130518 90510 131210 90536
rect 129904 90480 131210 90510
rect 131266 90480 131271 90536
rect 129904 90478 131271 90480
rect 129904 90450 130578 90478
rect 131205 90475 131271 90478
rect 131113 89994 131179 89997
rect 130518 89992 131179 89994
rect 130518 89966 131118 89992
rect 129904 89936 131118 89966
rect 131174 89936 131179 89992
rect 129904 89934 131179 89936
rect 129904 89906 130578 89934
rect 131113 89931 131179 89934
rect 186313 89994 186379 89997
rect 186313 89992 190164 89994
rect 186313 89936 186318 89992
rect 186374 89936 190164 89992
rect 186313 89934 190164 89936
rect 186313 89931 186379 89934
rect 411253 89722 411319 89725
rect 409860 89720 411319 89722
rect 409860 89664 411258 89720
rect 411314 89664 411319 89720
rect 409860 89662 411319 89664
rect 411253 89659 411319 89662
rect 437473 89586 437539 89589
rect 437473 89584 440066 89586
rect 437473 89528 437478 89584
rect 437534 89528 440066 89584
rect 437473 89526 440066 89528
rect 437473 89523 437539 89526
rect 132217 89450 132283 89453
rect 130518 89448 132283 89450
rect 130518 89422 132222 89448
rect 129904 89392 132222 89422
rect 132278 89392 132283 89448
rect 129904 89390 132283 89392
rect 129904 89362 130578 89390
rect 132217 89387 132283 89390
rect 440006 89148 440066 89526
rect 542353 89042 542419 89045
rect 539948 89040 542419 89042
rect 539948 88984 542358 89040
rect 542414 88984 542419 89040
rect 539948 88982 542419 88984
rect 542353 88979 542419 88982
rect 186313 88906 186379 88909
rect 186313 88904 190164 88906
rect 186313 88848 186318 88904
rect 186374 88848 190164 88904
rect 186313 88846 190164 88848
rect 186313 88843 186379 88846
rect 131297 88770 131363 88773
rect 130518 88768 131363 88770
rect 130518 88742 131302 88768
rect 129904 88712 131302 88742
rect 131358 88712 131363 88768
rect 129904 88710 131363 88712
rect 129904 88682 130578 88710
rect 131297 88707 131363 88710
rect 131205 88226 131271 88229
rect 130518 88224 131271 88226
rect 130518 88198 131210 88224
rect 129904 88168 131210 88198
rect 131266 88168 131271 88224
rect 129904 88166 131271 88168
rect 129904 88138 130578 88166
rect 131205 88163 131271 88166
rect 437473 87954 437539 87957
rect 437473 87952 440066 87954
rect 437473 87896 437478 87952
rect 437534 87896 440066 87952
rect 437473 87894 440066 87896
rect 437473 87891 437539 87894
rect 411253 87818 411319 87821
rect 409860 87816 411319 87818
rect 409860 87760 411258 87816
rect 411314 87760 411319 87816
rect 409860 87758 411319 87760
rect 411253 87755 411319 87758
rect 131113 87682 131179 87685
rect 130518 87680 131179 87682
rect 130518 87654 131118 87680
rect 129904 87624 131118 87654
rect 131174 87624 131179 87680
rect 129904 87622 131179 87624
rect 129904 87594 130578 87622
rect 131113 87619 131179 87622
rect 186313 87682 186379 87685
rect 186313 87680 190164 87682
rect 186313 87624 186318 87680
rect 186374 87624 190164 87680
rect 186313 87622 190164 87624
rect 186313 87619 186379 87622
rect 440006 87516 440066 87894
rect 131297 87002 131363 87005
rect 130518 87000 131363 87002
rect 130518 86974 131302 87000
rect 129904 86944 131302 86974
rect 131358 86944 131363 87000
rect 129904 86942 131363 86944
rect 129904 86914 130578 86942
rect 131297 86939 131363 86942
rect 131205 86458 131271 86461
rect 130518 86456 131271 86458
rect 130518 86430 131210 86456
rect 129904 86400 131210 86430
rect 131266 86400 131271 86456
rect 129904 86398 131271 86400
rect 129904 86370 130578 86398
rect 131205 86395 131271 86398
rect 186313 86458 186379 86461
rect 437473 86458 437539 86461
rect 186313 86456 190164 86458
rect 186313 86400 186318 86456
rect 186374 86400 190164 86456
rect 186313 86398 190164 86400
rect 437473 86456 440066 86458
rect 437473 86400 437478 86456
rect 437534 86400 440066 86456
rect 437473 86398 440066 86400
rect 186313 86395 186379 86398
rect 437473 86395 437539 86398
rect 131113 85914 131179 85917
rect 411253 85914 411319 85917
rect 130518 85912 131179 85914
rect 130518 85886 131118 85912
rect 129904 85856 131118 85886
rect 131174 85856 131179 85912
rect 129904 85854 131179 85856
rect 409860 85912 411319 85914
rect 409860 85856 411258 85912
rect 411314 85856 411319 85912
rect 440006 85884 440066 86398
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 409860 85854 411319 85856
rect 129904 85826 130578 85854
rect 131113 85851 131179 85854
rect 411253 85851 411319 85854
rect 132217 85370 132283 85373
rect 130518 85368 132283 85370
rect 130518 85342 132222 85368
rect 129904 85312 132222 85342
rect 132278 85312 132283 85368
rect 129904 85310 132283 85312
rect 129904 85282 130578 85310
rect 132217 85307 132283 85310
rect 187049 85370 187115 85373
rect 187049 85368 190164 85370
rect 187049 85312 187054 85368
rect 187110 85312 190164 85368
rect 187049 85310 190164 85312
rect 187049 85307 187115 85310
rect 437473 84826 437539 84829
rect 437473 84824 440066 84826
rect -960 84540 480 84780
rect 437473 84768 437478 84824
rect 437534 84768 440066 84824
rect 437473 84766 440066 84768
rect 437473 84763 437539 84766
rect 131113 84690 131179 84693
rect 130518 84688 131179 84690
rect 130518 84662 131118 84688
rect 129904 84632 131118 84662
rect 131174 84632 131179 84688
rect 129904 84630 131179 84632
rect 129904 84602 130578 84630
rect 131113 84627 131179 84630
rect 440006 84252 440066 84766
rect 132217 84146 132283 84149
rect 130518 84144 132283 84146
rect 130518 84118 132222 84144
rect 129904 84088 132222 84118
rect 132278 84088 132283 84144
rect 129904 84086 132283 84088
rect 129904 84058 130578 84086
rect 132217 84083 132283 84086
rect 186405 84146 186471 84149
rect 186405 84144 190164 84146
rect 186405 84088 186410 84144
rect 186466 84088 190164 84144
rect 186405 84086 190164 84088
rect 186405 84083 186471 84086
rect 411253 84010 411319 84013
rect 409860 84008 411319 84010
rect 409860 83952 411258 84008
rect 411314 83952 411319 84008
rect 409860 83950 411319 83952
rect 411253 83947 411319 83950
rect 131205 83602 131271 83605
rect 130518 83600 131271 83602
rect 130518 83574 131210 83600
rect 129904 83544 131210 83574
rect 131266 83544 131271 83600
rect 129904 83542 131271 83544
rect 129904 83514 130578 83542
rect 131205 83539 131271 83542
rect 186313 83058 186379 83061
rect 186313 83056 190164 83058
rect 186313 83000 186318 83056
rect 186374 83000 190164 83056
rect 186313 82998 190164 83000
rect 186313 82995 186379 82998
rect 131113 82922 131179 82925
rect 130518 82920 131179 82922
rect 130518 82894 131118 82920
rect 129904 82864 131118 82894
rect 131174 82864 131179 82920
rect 129904 82862 131179 82864
rect 129904 82834 130578 82862
rect 131113 82859 131179 82862
rect 437473 82786 437539 82789
rect 437473 82784 440066 82786
rect 437473 82728 437478 82784
rect 437534 82728 440066 82784
rect 437473 82726 440066 82728
rect 437473 82723 437539 82726
rect 440006 82484 440066 82726
rect 131573 82378 131639 82381
rect 130518 82376 131639 82378
rect 130518 82350 131578 82376
rect 129904 82320 131578 82350
rect 131634 82320 131639 82376
rect 129904 82318 131639 82320
rect 129904 82290 130578 82318
rect 131573 82315 131639 82318
rect 412449 82106 412515 82109
rect 409860 82104 412515 82106
rect 409860 82048 412454 82104
rect 412510 82048 412515 82104
rect 409860 82046 412515 82048
rect 412449 82043 412515 82046
rect 131205 81834 131271 81837
rect 130518 81832 131271 81834
rect 130518 81806 131210 81832
rect 129904 81776 131210 81806
rect 131266 81776 131271 81832
rect 129904 81774 131271 81776
rect 129904 81746 130578 81774
rect 131205 81771 131271 81774
rect 187141 81834 187207 81837
rect 187141 81832 190164 81834
rect 187141 81776 187146 81832
rect 187202 81776 190164 81832
rect 187141 81774 190164 81776
rect 187141 81771 187207 81774
rect 437473 81290 437539 81293
rect 437473 81288 440066 81290
rect 437473 81232 437478 81288
rect 437534 81232 440066 81288
rect 437473 81230 440066 81232
rect 437473 81227 437539 81230
rect 132217 81154 132283 81157
rect 130518 81152 132283 81154
rect 130518 81126 132222 81152
rect 129904 81096 132222 81126
rect 132278 81096 132283 81152
rect 129904 81094 132283 81096
rect 129904 81066 130578 81094
rect 132217 81091 132283 81094
rect 440006 80852 440066 81230
rect 186313 80746 186379 80749
rect 186313 80744 190164 80746
rect 186313 80688 186318 80744
rect 186374 80688 190164 80744
rect 186313 80686 190164 80688
rect 186313 80683 186379 80686
rect 131205 80610 131271 80613
rect 130518 80608 131271 80610
rect 130518 80582 131210 80608
rect 129904 80552 131210 80582
rect 131266 80552 131271 80608
rect 129904 80550 131271 80552
rect 129904 80522 130578 80550
rect 131205 80547 131271 80550
rect 411253 80202 411319 80205
rect 409860 80200 411319 80202
rect 409860 80144 411258 80200
rect 411314 80144 411319 80200
rect 409860 80142 411319 80144
rect 411253 80139 411319 80142
rect 131205 80066 131271 80069
rect 542445 80066 542511 80069
rect 130518 80064 131271 80066
rect 130518 80038 131210 80064
rect 129904 80008 131210 80038
rect 131266 80008 131271 80064
rect 129904 80006 131271 80008
rect 539948 80064 542511 80066
rect 539948 80008 542450 80064
rect 542506 80008 542511 80064
rect 539948 80006 542511 80008
rect 129904 79978 130578 80006
rect 131205 80003 131271 80006
rect 542445 80003 542511 80006
rect 437473 79658 437539 79661
rect 437473 79656 440066 79658
rect 437473 79600 437478 79656
rect 437534 79600 440066 79656
rect 437473 79598 440066 79600
rect 437473 79595 437539 79598
rect 131113 79522 131179 79525
rect 130518 79520 131179 79522
rect 130518 79494 131118 79520
rect 129904 79464 131118 79494
rect 131174 79464 131179 79520
rect 129904 79462 131179 79464
rect 129904 79434 130578 79462
rect 131113 79459 131179 79462
rect 186313 79522 186379 79525
rect 186313 79520 190164 79522
rect 186313 79464 186318 79520
rect 186374 79464 190164 79520
rect 186313 79462 190164 79464
rect 186313 79459 186379 79462
rect 440006 79220 440066 79598
rect 131205 78842 131271 78845
rect 130518 78840 131271 78842
rect 130518 78814 131210 78840
rect 129904 78784 131210 78814
rect 131266 78784 131271 78840
rect 129904 78782 131271 78784
rect 129904 78754 130578 78782
rect 131205 78779 131271 78782
rect 131205 78298 131271 78301
rect 130518 78296 131271 78298
rect 130518 78270 131210 78296
rect 129904 78240 131210 78270
rect 131266 78240 131271 78296
rect 129904 78238 131271 78240
rect 129904 78210 130578 78238
rect 131205 78235 131271 78238
rect 187417 78298 187483 78301
rect 411253 78298 411319 78301
rect 187417 78296 190164 78298
rect 187417 78240 187422 78296
rect 187478 78240 190164 78296
rect 187417 78238 190164 78240
rect 409860 78296 411319 78298
rect 409860 78240 411258 78296
rect 411314 78240 411319 78296
rect 409860 78238 411319 78240
rect 187417 78235 187483 78238
rect 411253 78235 411319 78238
rect 437473 78162 437539 78165
rect 437473 78160 440066 78162
rect 437473 78104 437478 78160
rect 437534 78104 440066 78160
rect 437473 78102 440066 78104
rect 437473 78099 437539 78102
rect 131113 77754 131179 77757
rect 130518 77752 131179 77754
rect 130518 77726 131118 77752
rect 129904 77696 131118 77726
rect 131174 77696 131179 77752
rect 129904 77694 131179 77696
rect 129904 77666 130578 77694
rect 131113 77691 131179 77694
rect 440006 77588 440066 78102
rect 186405 77210 186471 77213
rect 186405 77208 190164 77210
rect 186405 77152 186410 77208
rect 186466 77152 190164 77208
rect 186405 77150 190164 77152
rect 186405 77147 186471 77150
rect 131297 77074 131363 77077
rect 130518 77072 131363 77074
rect 130518 77046 131302 77072
rect 129904 77016 131302 77046
rect 131358 77016 131363 77072
rect 129904 77014 131363 77016
rect 129904 76986 130578 77014
rect 131297 77011 131363 77014
rect 131205 76530 131271 76533
rect 130518 76528 131271 76530
rect 130518 76502 131210 76528
rect 129904 76472 131210 76502
rect 131266 76472 131271 76528
rect 129904 76470 131271 76472
rect 129904 76442 130578 76470
rect 131205 76467 131271 76470
rect 411253 76394 411319 76397
rect 409860 76392 411319 76394
rect 409860 76336 411258 76392
rect 411314 76336 411319 76392
rect 409860 76334 411319 76336
rect 411253 76331 411319 76334
rect 131113 75986 131179 75989
rect 130518 75984 131179 75986
rect 130518 75958 131118 75984
rect 129904 75928 131118 75958
rect 131174 75928 131179 75984
rect 129904 75926 131179 75928
rect 129904 75898 130578 75926
rect 131113 75923 131179 75926
rect 186313 75986 186379 75989
rect 186313 75984 190164 75986
rect 186313 75928 186318 75984
rect 186374 75928 190164 75984
rect 186313 75926 190164 75928
rect 186313 75923 186379 75926
rect 437473 75714 437539 75717
rect 440006 75714 440066 75820
rect 437473 75712 440066 75714
rect 437473 75656 437478 75712
rect 437534 75656 440066 75712
rect 437473 75654 440066 75656
rect 437473 75651 437539 75654
rect 131205 75306 131271 75309
rect 130518 75304 131271 75306
rect 130518 75278 131210 75304
rect 129904 75248 131210 75278
rect 131266 75248 131271 75304
rect 129904 75246 131271 75248
rect 129904 75218 130578 75246
rect 131205 75243 131271 75246
rect 187233 74898 187299 74901
rect 187233 74896 190164 74898
rect 187233 74840 187238 74896
rect 187294 74840 190164 74896
rect 187233 74838 190164 74840
rect 187233 74835 187299 74838
rect 131113 74762 131179 74765
rect 130518 74760 131179 74762
rect 130518 74734 131118 74760
rect 129904 74704 131118 74734
rect 131174 74704 131179 74760
rect 129904 74702 131179 74704
rect 129904 74674 130578 74702
rect 131113 74699 131179 74702
rect 411253 74490 411319 74493
rect 409860 74488 411319 74490
rect 409860 74432 411258 74488
rect 411314 74432 411319 74488
rect 409860 74430 411319 74432
rect 411253 74427 411319 74430
rect 437473 74354 437539 74357
rect 437473 74352 440066 74354
rect 437473 74296 437478 74352
rect 437534 74296 440066 74352
rect 437473 74294 440066 74296
rect 437473 74291 437539 74294
rect 131205 74218 131271 74221
rect 130518 74216 131271 74218
rect 130518 74190 131210 74216
rect 129904 74160 131210 74190
rect 131266 74160 131271 74216
rect 440006 74188 440066 74294
rect 129904 74158 131271 74160
rect 129904 74130 130578 74158
rect 131205 74155 131271 74158
rect 131113 73674 131179 73677
rect 130518 73672 131179 73674
rect 130518 73646 131118 73672
rect 129904 73616 131118 73646
rect 131174 73616 131179 73672
rect 129904 73614 131179 73616
rect 129904 73586 130578 73614
rect 131113 73611 131179 73614
rect 186313 73674 186379 73677
rect 186313 73672 190164 73674
rect 186313 73616 186318 73672
rect 186374 73616 190164 73672
rect 186313 73614 190164 73616
rect 186313 73611 186379 73614
rect 131205 72994 131271 72997
rect 130518 72992 131271 72994
rect 130518 72966 131210 72992
rect 129904 72936 131210 72966
rect 131266 72936 131271 72992
rect 129904 72934 131271 72936
rect 129904 72906 130578 72934
rect 131205 72931 131271 72934
rect 437473 72858 437539 72861
rect 437473 72856 440066 72858
rect 437473 72800 437478 72856
rect 437534 72800 440066 72856
rect 583520 72844 584960 73084
rect 437473 72798 440066 72800
rect 437473 72795 437539 72798
rect 186313 72586 186379 72589
rect 411253 72586 411319 72589
rect 186313 72584 190164 72586
rect 186313 72528 186318 72584
rect 186374 72528 190164 72584
rect 186313 72526 190164 72528
rect 409860 72584 411319 72586
rect 409860 72528 411258 72584
rect 411314 72528 411319 72584
rect 440006 72556 440066 72798
rect 409860 72526 411319 72528
rect 186313 72523 186379 72526
rect 411253 72523 411319 72526
rect 131113 72450 131179 72453
rect 130518 72448 131179 72450
rect 130518 72422 131118 72448
rect 129904 72392 131118 72422
rect 131174 72392 131179 72448
rect 129904 72390 131179 72392
rect 129904 72362 130578 72390
rect 131113 72387 131179 72390
rect 132493 71906 132559 71909
rect 130518 71904 132559 71906
rect 130518 71878 132498 71904
rect 129904 71848 132498 71878
rect 132554 71848 132559 71904
rect 129904 71846 132559 71848
rect 129904 71818 130578 71846
rect 132493 71843 132559 71846
rect -960 71484 480 71724
rect 186313 71362 186379 71365
rect 437473 71362 437539 71365
rect 186313 71360 190164 71362
rect 186313 71304 186318 71360
rect 186374 71304 190164 71360
rect 186313 71302 190164 71304
rect 437473 71360 440066 71362
rect 437473 71304 437478 71360
rect 437534 71304 440066 71360
rect 437473 71302 440066 71304
rect 186313 71299 186379 71302
rect 437473 71299 437539 71302
rect 131205 71226 131271 71229
rect 130518 71224 131271 71226
rect 130518 71198 131210 71224
rect 129904 71168 131210 71198
rect 131266 71168 131271 71224
rect 129904 71166 131271 71168
rect 129904 71138 130578 71166
rect 131205 71163 131271 71166
rect 440006 70924 440066 71302
rect 542537 70954 542603 70957
rect 539948 70952 542603 70954
rect 539948 70896 542542 70952
rect 542598 70896 542603 70952
rect 539948 70894 542603 70896
rect 542537 70891 542603 70894
rect 131113 70682 131179 70685
rect 412357 70682 412423 70685
rect 130518 70680 131179 70682
rect 130518 70654 131118 70680
rect 129904 70624 131118 70654
rect 131174 70624 131179 70680
rect 129904 70622 131179 70624
rect 409860 70680 412423 70682
rect 409860 70624 412362 70680
rect 412418 70624 412423 70680
rect 409860 70622 412423 70624
rect 129904 70594 130578 70622
rect 131113 70619 131179 70622
rect 412357 70619 412423 70622
rect 186405 70274 186471 70277
rect 186405 70272 190164 70274
rect 186405 70216 186410 70272
rect 186466 70216 190164 70272
rect 186405 70214 190164 70216
rect 186405 70211 186471 70214
rect 131205 70138 131271 70141
rect 130518 70136 131271 70138
rect 130518 70110 131210 70136
rect 129904 70080 131210 70110
rect 131266 70080 131271 70136
rect 129904 70078 131271 70080
rect 129904 70050 130578 70078
rect 131205 70075 131271 70078
rect 437473 69730 437539 69733
rect 437473 69728 440066 69730
rect 437473 69672 437478 69728
rect 437534 69672 440066 69728
rect 437473 69670 440066 69672
rect 437473 69667 437539 69670
rect 131113 69458 131179 69461
rect 130518 69456 131179 69458
rect 130518 69430 131118 69456
rect 129904 69400 131118 69430
rect 131174 69400 131179 69456
rect 129904 69398 131179 69400
rect 129904 69370 130578 69398
rect 131113 69395 131179 69398
rect 440006 69156 440066 69670
rect 186313 69050 186379 69053
rect 186313 69048 190164 69050
rect 186313 68992 186318 69048
rect 186374 68992 190164 69048
rect 186313 68990 190164 68992
rect 186313 68987 186379 68990
rect 131113 68914 131179 68917
rect 130518 68912 131179 68914
rect 130518 68886 131118 68912
rect 129904 68856 131118 68886
rect 131174 68856 131179 68912
rect 129904 68854 131179 68856
rect 129904 68826 130578 68854
rect 131113 68851 131179 68854
rect 411345 68778 411411 68781
rect 409860 68776 411411 68778
rect 409860 68720 411350 68776
rect 411406 68720 411411 68776
rect 409860 68718 411411 68720
rect 411345 68715 411411 68718
rect 131205 68370 131271 68373
rect 130518 68368 131271 68370
rect 130518 68342 131210 68368
rect 129904 68312 131210 68342
rect 131266 68312 131271 68368
rect 129904 68310 131271 68312
rect 129904 68282 130578 68310
rect 131205 68307 131271 68310
rect 131297 67826 131363 67829
rect 130518 67824 131363 67826
rect 130518 67798 131302 67824
rect 129904 67768 131302 67798
rect 131358 67768 131363 67824
rect 129904 67766 131363 67768
rect 129904 67738 130578 67766
rect 131297 67763 131363 67766
rect 186313 67826 186379 67829
rect 186313 67824 190164 67826
rect 186313 67768 186318 67824
rect 186374 67768 190164 67824
rect 186313 67766 190164 67768
rect 186313 67763 186379 67766
rect 437473 67418 437539 67421
rect 440006 67418 440066 67524
rect 437473 67416 440066 67418
rect 437473 67360 437478 67416
rect 437534 67360 440066 67416
rect 437473 67358 440066 67360
rect 437473 67355 437539 67358
rect 131205 67146 131271 67149
rect 130518 67144 131271 67146
rect 130518 67118 131210 67144
rect 129904 67088 131210 67118
rect 131266 67088 131271 67144
rect 129904 67086 131271 67088
rect 129904 67058 130578 67086
rect 131205 67083 131271 67086
rect 411253 67010 411319 67013
rect 409860 67008 411319 67010
rect 409860 66952 411258 67008
rect 411314 66952 411319 67008
rect 409860 66950 411319 66952
rect 411253 66947 411319 66950
rect 186313 66738 186379 66741
rect 186313 66736 190164 66738
rect 186313 66680 186318 66736
rect 186374 66680 190164 66736
rect 186313 66678 190164 66680
rect 186313 66675 186379 66678
rect 131113 66602 131179 66605
rect 130518 66600 131179 66602
rect 130518 66574 131118 66600
rect 129904 66544 131118 66574
rect 131174 66544 131179 66600
rect 129904 66542 131179 66544
rect 129904 66514 130578 66542
rect 131113 66539 131179 66542
rect 437473 66194 437539 66197
rect 437473 66192 440066 66194
rect 437473 66136 437478 66192
rect 437534 66136 440066 66192
rect 437473 66134 440066 66136
rect 437473 66131 437539 66134
rect 131205 66058 131271 66061
rect 130518 66056 131271 66058
rect 130518 66030 131210 66056
rect 129904 66000 131210 66030
rect 131266 66000 131271 66056
rect 129904 65998 131271 66000
rect 129904 65970 130578 65998
rect 131205 65995 131271 65998
rect 440006 65892 440066 66134
rect 186313 65514 186379 65517
rect 186313 65512 190164 65514
rect 186313 65456 186318 65512
rect 186374 65456 190164 65512
rect 186313 65454 190164 65456
rect 186313 65451 186379 65454
rect 131113 65378 131179 65381
rect 130518 65376 131179 65378
rect 130518 65350 131118 65376
rect 129904 65320 131118 65350
rect 131174 65320 131179 65376
rect 129904 65318 131179 65320
rect 129904 65290 130578 65318
rect 131113 65315 131179 65318
rect 411253 65106 411319 65109
rect 409860 65104 411319 65106
rect 409860 65048 411258 65104
rect 411314 65048 411319 65104
rect 409860 65046 411319 65048
rect 411253 65043 411319 65046
rect 131205 64834 131271 64837
rect 130518 64832 131271 64834
rect 130518 64806 131210 64832
rect 129904 64776 131210 64806
rect 131266 64776 131271 64832
rect 129904 64774 131271 64776
rect 129904 64746 130578 64774
rect 131205 64771 131271 64774
rect 437473 64562 437539 64565
rect 437473 64560 440066 64562
rect 437473 64504 437478 64560
rect 437534 64504 440066 64560
rect 437473 64502 440066 64504
rect 437473 64499 437539 64502
rect 186313 64426 186379 64429
rect 186313 64424 190164 64426
rect 186313 64368 186318 64424
rect 186374 64368 190164 64424
rect 186313 64366 190164 64368
rect 186313 64363 186379 64366
rect 131849 64290 131915 64293
rect 130518 64288 131915 64290
rect 130518 64262 131854 64288
rect 129904 64232 131854 64262
rect 131910 64232 131915 64288
rect 440006 64260 440066 64502
rect 129904 64230 131915 64232
rect 129904 64202 130578 64230
rect 131849 64227 131915 64230
rect 131113 63746 131179 63749
rect 130518 63744 131179 63746
rect 130518 63718 131118 63744
rect 129904 63688 131118 63718
rect 131174 63688 131179 63744
rect 129904 63686 131179 63688
rect 129904 63658 130578 63686
rect 131113 63683 131179 63686
rect 186313 63202 186379 63205
rect 411253 63202 411319 63205
rect 186313 63200 190164 63202
rect 186313 63144 186318 63200
rect 186374 63144 190164 63200
rect 186313 63142 190164 63144
rect 409860 63200 411319 63202
rect 409860 63144 411258 63200
rect 411314 63144 411319 63200
rect 409860 63142 411319 63144
rect 186313 63139 186379 63142
rect 411253 63139 411319 63142
rect 132217 63066 132283 63069
rect 130518 63064 132283 63066
rect 130518 63038 132222 63064
rect 129904 63008 132222 63038
rect 132278 63008 132283 63064
rect 129904 63006 132283 63008
rect 129904 62978 130578 63006
rect 132217 63003 132283 63006
rect 438301 63066 438367 63069
rect 438301 63064 440066 63066
rect 438301 63008 438306 63064
rect 438362 63008 440066 63064
rect 438301 63006 440066 63008
rect 438301 63003 438367 63006
rect 131941 62522 132007 62525
rect 130518 62520 132007 62522
rect 130518 62494 131946 62520
rect 129904 62464 131946 62494
rect 132002 62464 132007 62520
rect 440006 62492 440066 63006
rect 129904 62462 132007 62464
rect 129904 62434 130578 62462
rect 131941 62459 132007 62462
rect 186405 62114 186471 62117
rect 186405 62112 190164 62114
rect 186405 62056 186410 62112
rect 186466 62056 190164 62112
rect 186405 62054 190164 62056
rect 186405 62051 186471 62054
rect 131205 61978 131271 61981
rect 130518 61976 131271 61978
rect 130518 61950 131210 61976
rect 129904 61920 131210 61950
rect 131266 61920 131271 61976
rect 129904 61918 131271 61920
rect 129904 61890 130578 61918
rect 131205 61915 131271 61918
rect 542629 61842 542695 61845
rect 539948 61840 542695 61842
rect 539948 61784 542634 61840
rect 542690 61784 542695 61840
rect 539948 61782 542695 61784
rect 542629 61779 542695 61782
rect 437473 61434 437539 61437
rect 437473 61432 440066 61434
rect 437473 61376 437478 61432
rect 437534 61376 440066 61432
rect 437473 61374 440066 61376
rect 437473 61371 437539 61374
rect 132125 61298 132191 61301
rect 411253 61298 411319 61301
rect 130518 61296 132191 61298
rect 130518 61270 132130 61296
rect 129904 61240 132130 61270
rect 132186 61240 132191 61296
rect 129904 61238 132191 61240
rect 409860 61296 411319 61298
rect 409860 61240 411258 61296
rect 411314 61240 411319 61296
rect 409860 61238 411319 61240
rect 129904 61210 130578 61238
rect 132125 61235 132191 61238
rect 411253 61235 411319 61238
rect 186313 60890 186379 60893
rect 186313 60888 190164 60890
rect 186313 60832 186318 60888
rect 186374 60832 190164 60888
rect 440006 60860 440066 61374
rect 186313 60830 190164 60832
rect 186313 60827 186379 60830
rect 131113 60754 131179 60757
rect 130150 60752 131179 60754
rect 130150 60720 131118 60752
rect 129904 60696 131118 60720
rect 131174 60696 131179 60752
rect 129904 60694 131179 60696
rect 129904 60660 130210 60694
rect 131113 60691 131179 60694
rect 132217 60210 132283 60213
rect 130518 60208 132283 60210
rect 130518 60182 132222 60208
rect 129904 60152 132222 60182
rect 132278 60152 132283 60208
rect 129904 60150 132283 60152
rect 129904 60122 130578 60150
rect 132217 60147 132283 60150
rect 186313 59802 186379 59805
rect 186313 59800 190164 59802
rect 186313 59744 186318 59800
rect 186374 59744 190164 59800
rect 186313 59742 190164 59744
rect 186313 59739 186379 59742
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 131665 59530 131731 59533
rect 130518 59528 131731 59530
rect 130518 59502 131670 59528
rect 129904 59472 131670 59502
rect 131726 59472 131731 59528
rect 583520 59516 584960 59606
rect 129904 59470 131731 59472
rect 129904 59442 130578 59470
rect 131665 59467 131731 59470
rect 411345 59394 411411 59397
rect 409860 59392 411411 59394
rect 409860 59336 411350 59392
rect 411406 59336 411411 59392
rect 409860 59334 411411 59336
rect 411345 59331 411411 59334
rect 437473 59122 437539 59125
rect 440006 59122 440066 59228
rect 437473 59120 440066 59122
rect 437473 59064 437478 59120
rect 437534 59064 440066 59120
rect 437473 59062 440066 59064
rect 437473 59059 437539 59062
rect 132033 58986 132099 58989
rect 130518 58984 132099 58986
rect 130518 58958 132038 58984
rect 129904 58928 132038 58958
rect 132094 58928 132099 58984
rect 129904 58926 132099 58928
rect 129904 58898 130578 58926
rect 132033 58923 132099 58926
rect -960 58428 480 58668
rect 186313 58578 186379 58581
rect 186313 58576 190164 58578
rect 186313 58520 186318 58576
rect 186374 58520 190164 58576
rect 186313 58518 190164 58520
rect 186313 58515 186379 58518
rect 131297 58442 131363 58445
rect 130518 58440 131363 58442
rect 130518 58414 131302 58440
rect 129904 58384 131302 58414
rect 131358 58384 131363 58440
rect 129904 58382 131363 58384
rect 129904 58354 130578 58382
rect 131297 58379 131363 58382
rect 131205 57898 131271 57901
rect 130518 57896 131271 57898
rect 130518 57870 131210 57896
rect 129904 57840 131210 57870
rect 131266 57840 131271 57896
rect 129904 57838 131271 57840
rect 129904 57810 130578 57838
rect 131205 57835 131271 57838
rect 437473 57898 437539 57901
rect 437473 57896 440066 57898
rect 437473 57840 437478 57896
rect 437534 57840 440066 57896
rect 437473 57838 440066 57840
rect 437473 57835 437539 57838
rect 440006 57596 440066 57838
rect 411253 57490 411319 57493
rect 409860 57488 411319 57490
rect 409860 57432 411258 57488
rect 411314 57432 411319 57488
rect 409860 57430 411319 57432
rect 411253 57427 411319 57430
rect 186957 57354 187023 57357
rect 186957 57352 190164 57354
rect 186957 57296 186962 57352
rect 187018 57296 190164 57352
rect 186957 57294 190164 57296
rect 186957 57291 187023 57294
rect 131205 57218 131271 57221
rect 130518 57216 131271 57218
rect 130518 57190 131210 57216
rect 129904 57160 131210 57190
rect 131266 57160 131271 57216
rect 129904 57158 131271 57160
rect 129904 57130 130578 57158
rect 131205 57155 131271 57158
rect 131113 56674 131179 56677
rect 130518 56672 131179 56674
rect 130518 56646 131118 56672
rect 129904 56616 131118 56646
rect 131174 56616 131179 56672
rect 129904 56614 131179 56616
rect 129904 56586 130578 56614
rect 131113 56611 131179 56614
rect 437749 56402 437815 56405
rect 437749 56400 440066 56402
rect 437749 56344 437754 56400
rect 437810 56344 440066 56400
rect 437749 56342 440066 56344
rect 437749 56339 437815 56342
rect 186313 56266 186379 56269
rect 186313 56264 190164 56266
rect 186313 56208 186318 56264
rect 186374 56208 190164 56264
rect 186313 56206 190164 56208
rect 186313 56203 186379 56206
rect 132217 56130 132283 56133
rect 130518 56128 132283 56130
rect 130518 56102 132222 56128
rect 129904 56072 132222 56102
rect 132278 56072 132283 56128
rect 129904 56070 132283 56072
rect 129904 56042 130578 56070
rect 132217 56067 132283 56070
rect 440006 55828 440066 56342
rect 411253 55586 411319 55589
rect 409860 55584 411319 55586
rect 409860 55528 411258 55584
rect 411314 55528 411319 55584
rect 409860 55526 411319 55528
rect 411253 55523 411319 55526
rect 131205 55450 131271 55453
rect 130518 55448 131271 55450
rect 130518 55422 131210 55448
rect 129904 55392 131210 55422
rect 131266 55392 131271 55448
rect 129904 55390 131271 55392
rect 129904 55362 130578 55390
rect 131205 55387 131271 55390
rect 186313 55042 186379 55045
rect 186313 55040 190164 55042
rect 186313 54984 186318 55040
rect 186374 54984 190164 55040
rect 186313 54982 190164 54984
rect 186313 54979 186379 54982
rect 131205 54906 131271 54909
rect 130518 54904 131271 54906
rect 130518 54878 131210 54904
rect 129904 54848 131210 54878
rect 131266 54848 131271 54904
rect 129904 54846 131271 54848
rect 129904 54818 130578 54846
rect 131205 54843 131271 54846
rect 437473 54770 437539 54773
rect 437473 54768 440066 54770
rect 437473 54712 437478 54768
rect 437534 54712 440066 54768
rect 437473 54710 440066 54712
rect 437473 54707 437539 54710
rect 132493 54362 132559 54365
rect 130518 54360 132559 54362
rect 130518 54334 132498 54360
rect 129904 54304 132498 54334
rect 132554 54304 132559 54360
rect 129904 54302 132559 54304
rect 129904 54274 130578 54302
rect 132493 54299 132559 54302
rect 440006 54196 440066 54710
rect 187049 53954 187115 53957
rect 187049 53952 190164 53954
rect 187049 53896 187054 53952
rect 187110 53896 190164 53952
rect 187049 53894 190164 53896
rect 187049 53891 187115 53894
rect 131297 53682 131363 53685
rect 412265 53682 412331 53685
rect 130518 53680 131363 53682
rect 130518 53654 131302 53680
rect 129904 53624 131302 53654
rect 131358 53624 131363 53680
rect 129904 53622 131363 53624
rect 409860 53680 412331 53682
rect 409860 53624 412270 53680
rect 412326 53624 412331 53680
rect 409860 53622 412331 53624
rect 129904 53594 130578 53622
rect 131297 53619 131363 53622
rect 412265 53619 412331 53622
rect 131205 53138 131271 53141
rect 130518 53136 131271 53138
rect 130518 53110 131210 53136
rect 129904 53080 131210 53110
rect 131266 53080 131271 53136
rect 129904 53078 131271 53080
rect 129904 53050 130578 53078
rect 131205 53075 131271 53078
rect 437473 53138 437539 53141
rect 437473 53136 440066 53138
rect 437473 53080 437478 53136
rect 437534 53080 440066 53136
rect 437473 53078 440066 53080
rect 437473 53075 437539 53078
rect 186313 52730 186379 52733
rect 186313 52728 190164 52730
rect 186313 52672 186318 52728
rect 186374 52672 190164 52728
rect 186313 52670 190164 52672
rect 186313 52667 186379 52670
rect 131113 52594 131179 52597
rect 130518 52592 131179 52594
rect 130518 52566 131118 52592
rect 129904 52536 131118 52566
rect 131174 52536 131179 52592
rect 440006 52564 440066 53078
rect 542721 52730 542787 52733
rect 539948 52728 542787 52730
rect 539948 52672 542726 52728
rect 542782 52672 542787 52728
rect 539948 52670 542787 52672
rect 542721 52667 542787 52670
rect 129904 52534 131179 52536
rect 129904 52506 130578 52534
rect 131113 52531 131179 52534
rect 132309 52050 132375 52053
rect 130518 52048 132375 52050
rect 130518 52022 132314 52048
rect 129904 51992 132314 52022
rect 132370 51992 132375 52048
rect 129904 51990 132375 51992
rect 129904 51962 130578 51990
rect 132309 51987 132375 51990
rect 412357 51778 412423 51781
rect 409860 51776 412423 51778
rect 409860 51720 412362 51776
rect 412418 51720 412423 51776
rect 409860 51718 412423 51720
rect 412357 51715 412423 51718
rect 186313 51642 186379 51645
rect 186313 51640 190164 51642
rect 186313 51584 186318 51640
rect 186374 51584 190164 51640
rect 186313 51582 190164 51584
rect 186313 51579 186379 51582
rect 131205 51370 131271 51373
rect 130518 51368 131271 51370
rect 130518 51342 131210 51368
rect 129904 51312 131210 51342
rect 131266 51312 131271 51368
rect 129904 51310 131271 51312
rect 129904 51282 130578 51310
rect 131205 51307 131271 51310
rect 131205 50826 131271 50829
rect 130518 50824 131271 50826
rect 130518 50798 131210 50824
rect 129904 50768 131210 50798
rect 131266 50768 131271 50824
rect 129904 50766 131271 50768
rect 129904 50738 130578 50766
rect 131205 50763 131271 50766
rect 436829 50826 436895 50829
rect 440006 50826 440066 50932
rect 436829 50824 440066 50826
rect 436829 50768 436834 50824
rect 436890 50768 440066 50824
rect 436829 50766 440066 50768
rect 436829 50763 436895 50766
rect 187141 50418 187207 50421
rect 187141 50416 190164 50418
rect 187141 50360 187146 50416
rect 187202 50360 190164 50416
rect 187141 50358 190164 50360
rect 187141 50355 187207 50358
rect 131113 50282 131179 50285
rect 130518 50280 131179 50282
rect 130518 50254 131118 50280
rect 129904 50224 131118 50254
rect 131174 50224 131179 50280
rect 129904 50222 131179 50224
rect 129904 50194 130578 50222
rect 131113 50219 131179 50222
rect 411253 49874 411319 49877
rect 409860 49872 411319 49874
rect 409860 49816 411258 49872
rect 411314 49816 411319 49872
rect 409860 49814 411319 49816
rect 411253 49811 411319 49814
rect 131297 49602 131363 49605
rect 130518 49600 131363 49602
rect 130518 49574 131302 49600
rect 129904 49544 131302 49574
rect 131358 49544 131363 49600
rect 129904 49542 131363 49544
rect 129904 49514 130578 49542
rect 131297 49539 131363 49542
rect 437473 49602 437539 49605
rect 437473 49600 440066 49602
rect 437473 49544 437478 49600
rect 437534 49544 440066 49600
rect 437473 49542 440066 49544
rect 437473 49539 437539 49542
rect 186313 49194 186379 49197
rect 186313 49192 190164 49194
rect 186313 49136 186318 49192
rect 186374 49136 190164 49192
rect 440006 49164 440066 49542
rect 186313 49134 190164 49136
rect 186313 49131 186379 49134
rect 131205 49058 131271 49061
rect 130518 49056 131271 49058
rect 130518 49030 131210 49056
rect 129904 49000 131210 49030
rect 131266 49000 131271 49056
rect 129904 48998 131271 49000
rect 129904 48970 130578 48998
rect 131205 48995 131271 48998
rect 131113 48514 131179 48517
rect 130518 48512 131179 48514
rect 130518 48486 131118 48512
rect 129904 48456 131118 48486
rect 131174 48456 131179 48512
rect 129904 48454 131179 48456
rect 129904 48426 130578 48454
rect 131113 48451 131179 48454
rect 186313 48106 186379 48109
rect 186313 48104 190164 48106
rect 186313 48048 186318 48104
rect 186374 48048 190164 48104
rect 186313 48046 190164 48048
rect 186313 48043 186379 48046
rect 411253 47970 411319 47973
rect 409860 47968 411319 47970
rect 409860 47912 411258 47968
rect 411314 47912 411319 47968
rect 409860 47910 411319 47912
rect 411253 47907 411319 47910
rect 437473 47970 437539 47973
rect 437473 47968 440066 47970
rect 437473 47912 437478 47968
rect 437534 47912 440066 47968
rect 437473 47910 440066 47912
rect 437473 47907 437539 47910
rect 131941 47834 132007 47837
rect 130518 47832 132007 47834
rect 130518 47806 131946 47832
rect 129904 47776 131946 47806
rect 132002 47776 132007 47832
rect 129904 47774 132007 47776
rect 129904 47746 130578 47774
rect 131941 47771 132007 47774
rect 440006 47532 440066 47910
rect 131205 47290 131271 47293
rect 130518 47288 131271 47290
rect 130518 47262 131210 47288
rect 129904 47232 131210 47262
rect 131266 47232 131271 47288
rect 129904 47230 131271 47232
rect 129904 47202 130578 47230
rect 131205 47227 131271 47230
rect 187417 46882 187483 46885
rect 187417 46880 190164 46882
rect 187417 46824 187422 46880
rect 187478 46824 190164 46880
rect 187417 46822 190164 46824
rect 187417 46819 187483 46822
rect 131205 46746 131271 46749
rect 130518 46744 131271 46746
rect 130518 46718 131210 46744
rect 129904 46688 131210 46718
rect 131266 46688 131271 46744
rect 129904 46686 131271 46688
rect 129904 46658 130578 46686
rect 131205 46683 131271 46686
rect 437473 46474 437539 46477
rect 437473 46472 440066 46474
rect 437473 46416 437478 46472
rect 437534 46416 440066 46472
rect 437473 46414 440066 46416
rect 437473 46411 437539 46414
rect 131113 46202 131179 46205
rect 130518 46200 131179 46202
rect 130518 46174 131118 46200
rect 129904 46144 131118 46174
rect 131174 46144 131179 46200
rect 129904 46142 131179 46144
rect 129904 46114 130578 46142
rect 131113 46139 131179 46142
rect 411253 46066 411319 46069
rect 409860 46064 411319 46066
rect 409860 46008 411258 46064
rect 411314 46008 411319 46064
rect 409860 46006 411319 46008
rect 411253 46003 411319 46006
rect 440006 45900 440066 46414
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect 187233 45794 187299 45797
rect 187233 45792 190164 45794
rect 187233 45736 187238 45792
rect 187294 45736 190164 45792
rect 187233 45734 190164 45736
rect 187233 45731 187299 45734
rect -960 45372 480 45612
rect 129968 45394 130578 45454
rect 130518 45386 130578 45394
rect 131205 45386 131271 45389
rect 130518 45384 131271 45386
rect 130518 45328 131210 45384
rect 131266 45328 131271 45384
rect 130518 45326 131271 45328
rect 131205 45323 131271 45326
rect 131113 44978 131179 44981
rect 130518 44976 131179 44978
rect 130518 44950 131118 44976
rect 129904 44920 131118 44950
rect 131174 44920 131179 44976
rect 129904 44918 131179 44920
rect 129904 44890 130578 44918
rect 131113 44915 131179 44918
rect 437473 44842 437539 44845
rect 437473 44840 440066 44842
rect 437473 44784 437478 44840
rect 437534 44784 440066 44840
rect 437473 44782 440066 44784
rect 437473 44779 437539 44782
rect 186313 44570 186379 44573
rect 186313 44568 190164 44570
rect 186313 44512 186318 44568
rect 186374 44512 190164 44568
rect 186313 44510 190164 44512
rect 186313 44507 186379 44510
rect 131297 44434 131363 44437
rect 130518 44432 131363 44434
rect 130518 44406 131302 44432
rect 129904 44376 131302 44406
rect 131358 44376 131363 44432
rect 129904 44374 131363 44376
rect 129904 44346 130578 44374
rect 131297 44371 131363 44374
rect 440006 44268 440066 44782
rect 411805 44162 411871 44165
rect 409860 44160 411871 44162
rect 409860 44104 411810 44160
rect 411866 44104 411871 44160
rect 409860 44102 411871 44104
rect 411805 44099 411871 44102
rect 131205 43754 131271 43757
rect 130518 43752 131271 43754
rect 130518 43726 131210 43752
rect 129904 43696 131210 43726
rect 131266 43696 131271 43752
rect 129904 43694 131271 43696
rect 129904 43666 130578 43694
rect 131205 43691 131271 43694
rect 542997 43618 543063 43621
rect 539948 43616 543063 43618
rect 539948 43560 543002 43616
rect 543058 43560 543063 43616
rect 539948 43558 543063 43560
rect 542997 43555 543063 43558
rect 186313 43482 186379 43485
rect 186313 43480 190164 43482
rect 186313 43424 186318 43480
rect 186374 43424 190164 43480
rect 186313 43422 190164 43424
rect 186313 43419 186379 43422
rect 131113 43210 131179 43213
rect 130518 43208 131179 43210
rect 130518 43182 131118 43208
rect 129904 43152 131118 43182
rect 131174 43152 131179 43208
rect 129904 43150 131179 43152
rect 129904 43122 130578 43150
rect 131113 43147 131179 43150
rect 131205 42666 131271 42669
rect 130518 42664 131271 42666
rect 130518 42638 131210 42664
rect 129904 42608 131210 42638
rect 131266 42608 131271 42664
rect 129904 42606 131271 42608
rect 129904 42578 130578 42606
rect 131205 42603 131271 42606
rect 437473 42666 437539 42669
rect 437473 42664 440066 42666
rect 437473 42608 437478 42664
rect 437534 42608 440066 42664
rect 437473 42606 440066 42608
rect 437473 42603 437539 42606
rect 440006 42500 440066 42606
rect 186405 42258 186471 42261
rect 411253 42258 411319 42261
rect 186405 42256 190164 42258
rect 186405 42200 186410 42256
rect 186466 42200 190164 42256
rect 186405 42198 190164 42200
rect 409860 42256 411319 42258
rect 409860 42200 411258 42256
rect 411314 42200 411319 42256
rect 409860 42198 411319 42200
rect 186405 42195 186471 42198
rect 411253 42195 411319 42198
rect 131113 41986 131179 41989
rect 130518 41984 131179 41986
rect 130518 41958 131118 41984
rect 129904 41928 131118 41958
rect 131174 41928 131179 41984
rect 129904 41926 131179 41928
rect 129904 41898 130578 41926
rect 131113 41923 131179 41926
rect 131849 41442 131915 41445
rect 130150 41440 131915 41442
rect 130150 41408 131854 41440
rect 129904 41384 131854 41408
rect 131910 41384 131915 41440
rect 129904 41382 131915 41384
rect 129904 41348 130210 41382
rect 131849 41379 131915 41382
rect 437473 41306 437539 41309
rect 437473 41304 440066 41306
rect 437473 41248 437478 41304
rect 437534 41248 440066 41304
rect 437473 41246 440066 41248
rect 437473 41243 437539 41246
rect 186957 41170 187023 41173
rect 186957 41168 190164 41170
rect 186957 41112 186962 41168
rect 187018 41112 190164 41168
rect 186957 41110 190164 41112
rect 186957 41107 187023 41110
rect 131205 40898 131271 40901
rect 130518 40896 131271 40898
rect 130518 40870 131210 40896
rect 129904 40840 131210 40870
rect 131266 40840 131271 40896
rect 440006 40868 440066 41246
rect 129904 40838 131271 40840
rect 129904 40810 130578 40838
rect 131205 40835 131271 40838
rect 131113 40354 131179 40357
rect 411253 40354 411319 40357
rect 130518 40352 131179 40354
rect 130518 40326 131118 40352
rect 129904 40296 131118 40326
rect 131174 40296 131179 40352
rect 129904 40294 131179 40296
rect 409860 40352 411319 40354
rect 409860 40296 411258 40352
rect 411314 40296 411319 40352
rect 409860 40294 411319 40296
rect 129904 40266 130578 40294
rect 131113 40291 131179 40294
rect 411253 40291 411319 40294
rect 187049 39946 187115 39949
rect 187049 39944 190164 39946
rect 187049 39888 187054 39944
rect 187110 39888 190164 39944
rect 187049 39886 190164 39888
rect 187049 39883 187115 39886
rect 131941 39674 132007 39677
rect 130518 39672 132007 39674
rect 130518 39646 131946 39672
rect 129904 39616 131946 39646
rect 132002 39616 132007 39672
rect 129904 39614 132007 39616
rect 129904 39586 130578 39614
rect 131941 39611 132007 39614
rect 437473 39674 437539 39677
rect 437473 39672 440066 39674
rect 437473 39616 437478 39672
rect 437534 39616 440066 39672
rect 437473 39614 440066 39616
rect 437473 39611 437539 39614
rect 440006 39236 440066 39614
rect 132493 39130 132559 39133
rect 130518 39128 132559 39130
rect 130518 39102 132498 39128
rect 129904 39072 132498 39102
rect 132554 39072 132559 39128
rect 129904 39070 132559 39072
rect 129904 39042 130578 39070
rect 132493 39067 132559 39070
rect 186313 38722 186379 38725
rect 186313 38720 190164 38722
rect 186313 38664 186318 38720
rect 186374 38664 190164 38720
rect 186313 38662 190164 38664
rect 186313 38659 186379 38662
rect 131205 38586 131271 38589
rect 130518 38584 131271 38586
rect 130518 38558 131210 38584
rect 129904 38528 131210 38558
rect 131266 38528 131271 38584
rect 129904 38526 131271 38528
rect 129904 38498 130578 38526
rect 131205 38523 131271 38526
rect 411253 38450 411319 38453
rect 409860 38448 411319 38450
rect 409860 38392 411258 38448
rect 411314 38392 411319 38448
rect 409860 38390 411319 38392
rect 411253 38387 411319 38390
rect 437473 38178 437539 38181
rect 437473 38176 440066 38178
rect 437473 38120 437478 38176
rect 437534 38120 440066 38176
rect 437473 38118 440066 38120
rect 437473 38115 437539 38118
rect 131113 37906 131179 37909
rect 130518 37904 131179 37906
rect 130518 37878 131118 37904
rect 129904 37848 131118 37878
rect 131174 37848 131179 37904
rect 129904 37846 131179 37848
rect 129904 37818 130578 37846
rect 131113 37843 131179 37846
rect 186313 37634 186379 37637
rect 186313 37632 190164 37634
rect 186313 37576 186318 37632
rect 186374 37576 190164 37632
rect 440006 37604 440066 38118
rect 186313 37574 190164 37576
rect 186313 37571 186379 37574
rect 131481 37362 131547 37365
rect 130518 37360 131547 37362
rect 130518 37334 131486 37360
rect 129904 37304 131486 37334
rect 131542 37304 131547 37360
rect 129904 37302 131547 37304
rect 129904 37274 130578 37302
rect 131481 37299 131547 37302
rect 131297 36818 131363 36821
rect 130518 36816 131363 36818
rect 130518 36790 131302 36816
rect 129904 36760 131302 36790
rect 131358 36760 131363 36816
rect 129904 36758 131363 36760
rect 129904 36730 130578 36758
rect 131297 36755 131363 36758
rect 411253 36546 411319 36549
rect 409860 36544 411319 36546
rect 409860 36488 411258 36544
rect 411314 36488 411319 36544
rect 409860 36486 411319 36488
rect 411253 36483 411319 36486
rect 186313 36410 186379 36413
rect 186313 36408 190164 36410
rect 186313 36352 186318 36408
rect 186374 36352 190164 36408
rect 186313 36350 190164 36352
rect 186313 36347 186379 36350
rect 131205 36138 131271 36141
rect 130518 36136 131271 36138
rect 130518 36110 131210 36136
rect 129904 36080 131210 36110
rect 131266 36080 131271 36136
rect 129904 36078 131271 36080
rect 129904 36050 130578 36078
rect 131205 36075 131271 36078
rect 437473 35730 437539 35733
rect 440006 35730 440066 35836
rect 437473 35728 440066 35730
rect 437473 35672 437478 35728
rect 437534 35672 440066 35728
rect 437473 35670 440066 35672
rect 437473 35667 437539 35670
rect 131205 35594 131271 35597
rect 130518 35592 131271 35594
rect 130518 35566 131210 35592
rect 129904 35536 131210 35566
rect 131266 35536 131271 35592
rect 129904 35534 131271 35536
rect 129904 35506 130578 35534
rect 131205 35531 131271 35534
rect 186405 35322 186471 35325
rect 186405 35320 190164 35322
rect 186405 35264 186410 35320
rect 186466 35264 190164 35320
rect 186405 35262 190164 35264
rect 186405 35259 186471 35262
rect 131113 35050 131179 35053
rect 130518 35048 131179 35050
rect 130518 35022 131118 35048
rect 129904 34992 131118 35022
rect 131174 34992 131179 35048
rect 129904 34990 131179 34992
rect 129904 34962 130578 34990
rect 131113 34987 131179 34990
rect 411253 34642 411319 34645
rect 543089 34642 543155 34645
rect 409860 34640 411319 34642
rect 409860 34584 411258 34640
rect 411314 34584 411319 34640
rect 409860 34582 411319 34584
rect 539948 34640 543155 34642
rect 539948 34584 543094 34640
rect 543150 34584 543155 34640
rect 539948 34582 543155 34584
rect 411253 34579 411319 34582
rect 543089 34579 543155 34582
rect 131849 34506 131915 34509
rect 130518 34504 131915 34506
rect 130518 34478 131854 34504
rect 129904 34448 131854 34478
rect 131910 34448 131915 34504
rect 129904 34446 131915 34448
rect 129904 34418 130578 34446
rect 131849 34443 131915 34446
rect 437473 34370 437539 34373
rect 437473 34368 440066 34370
rect 437473 34312 437478 34368
rect 437534 34312 440066 34368
rect 437473 34310 440066 34312
rect 437473 34307 437539 34310
rect 440006 34204 440066 34310
rect 186313 34098 186379 34101
rect 186313 34096 190164 34098
rect 186313 34040 186318 34096
rect 186374 34040 190164 34096
rect 186313 34038 190164 34040
rect 186313 34035 186379 34038
rect 132125 33826 132191 33829
rect 130518 33824 132191 33826
rect 130518 33798 132130 33824
rect 129904 33768 132130 33798
rect 132186 33768 132191 33824
rect 129904 33766 132191 33768
rect 129904 33738 130578 33766
rect 132125 33763 132191 33766
rect 132217 33282 132283 33285
rect 130518 33280 132283 33282
rect 130518 33254 132222 33280
rect 129904 33224 132222 33254
rect 132278 33224 132283 33280
rect 129904 33222 132283 33224
rect 129904 33194 130578 33222
rect 132217 33219 132283 33222
rect 186405 33010 186471 33013
rect 437473 33010 437539 33013
rect 186405 33008 190164 33010
rect 186405 32952 186410 33008
rect 186466 32952 190164 33008
rect 186405 32950 190164 32952
rect 437473 33008 440066 33010
rect 437473 32952 437478 33008
rect 437534 32952 440066 33008
rect 583520 32996 584960 33236
rect 437473 32950 440066 32952
rect 186405 32947 186471 32950
rect 437473 32947 437539 32950
rect 131205 32738 131271 32741
rect 411253 32738 411319 32741
rect 130518 32736 131271 32738
rect 130518 32710 131210 32736
rect 129904 32680 131210 32710
rect 131266 32680 131271 32736
rect 129904 32678 131271 32680
rect 409860 32736 411319 32738
rect 409860 32680 411258 32736
rect 411314 32680 411319 32736
rect 409860 32678 411319 32680
rect 129904 32650 130578 32678
rect 131205 32675 131271 32678
rect 411253 32675 411319 32678
rect 440006 32572 440066 32950
rect -960 32316 480 32556
rect 131113 32058 131179 32061
rect 130518 32056 131179 32058
rect 130518 32030 131118 32056
rect 129904 32000 131118 32030
rect 131174 32000 131179 32056
rect 129904 31998 131179 32000
rect 129904 31970 130578 31998
rect 131113 31995 131179 31998
rect 186313 31786 186379 31789
rect 186313 31784 190164 31786
rect 186313 31728 186318 31784
rect 186374 31728 190164 31784
rect 186313 31726 190164 31728
rect 186313 31723 186379 31726
rect 131205 31514 131271 31517
rect 130518 31512 131271 31514
rect 130518 31486 131210 31512
rect 129904 31456 131210 31486
rect 131266 31456 131271 31512
rect 129904 31454 131271 31456
rect 129904 31426 130578 31454
rect 131205 31451 131271 31454
rect 437473 31242 437539 31245
rect 437473 31240 440066 31242
rect 437473 31184 437478 31240
rect 437534 31184 440066 31240
rect 437473 31182 440066 31184
rect 437473 31179 437539 31182
rect 131297 30970 131363 30973
rect 411253 30970 411319 30973
rect 130518 30968 131363 30970
rect 130518 30942 131302 30968
rect 129904 30912 131302 30942
rect 131358 30912 131363 30968
rect 129904 30910 131363 30912
rect 409860 30968 411319 30970
rect 409860 30912 411258 30968
rect 411314 30912 411319 30968
rect 440006 30940 440066 31182
rect 409860 30910 411319 30912
rect 129904 30882 130578 30910
rect 131297 30907 131363 30910
rect 411253 30907 411319 30910
rect 186313 30698 186379 30701
rect 186313 30696 190164 30698
rect 186313 30640 186318 30696
rect 186374 30640 190164 30696
rect 186313 30638 190164 30640
rect 186313 30635 186379 30638
rect 131113 30426 131179 30429
rect 130150 30424 131179 30426
rect 129782 30290 129842 30396
rect 130150 30368 131118 30424
rect 131174 30368 131179 30424
rect 130150 30366 131179 30368
rect 130150 30290 130210 30366
rect 131113 30363 131179 30366
rect 129782 30230 130210 30290
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19260 480 19500
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6340 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 583520 6476 584960 6566
<< via3 >>
rect 239654 299780 239718 299844
rect 243054 299704 243118 299708
rect 243054 299648 243082 299704
rect 243082 299648 243118 299704
rect 243054 299644 243118 299648
rect 55854 299568 55918 299572
rect 55854 299512 55862 299568
rect 55862 299512 55918 299568
rect 55854 299508 55918 299512
rect 67822 299568 67886 299572
rect 67822 299512 67878 299568
rect 67878 299512 67886 299568
rect 67822 299508 67886 299512
rect 229140 298344 229204 298348
rect 229140 298288 229154 298344
rect 229154 298288 229204 298344
rect 229140 298284 229204 298288
rect 73660 298148 73724 298212
rect 77892 298148 77956 298212
rect 81756 298148 81820 298212
rect 85436 298148 85500 298212
rect 91876 298148 91940 298212
rect 95556 298148 95620 298212
rect 95924 298148 95988 298212
rect 99420 298148 99484 298212
rect 102916 298148 102980 298212
rect 103284 298148 103348 298212
rect 225460 298148 225524 298212
rect 257844 298148 257908 298212
rect 261524 298148 261588 298212
rect 261892 298148 261956 298212
rect 265204 298148 265268 298212
rect 271828 298148 271892 298212
rect 275508 298148 275572 298212
rect 65564 298012 65628 298076
rect 66668 298012 66732 298076
rect 69244 298072 69308 298076
rect 69244 298016 69294 298072
rect 69294 298016 69308 298072
rect 69244 298012 69308 298016
rect 70164 298072 70228 298076
rect 70164 298016 70214 298072
rect 70214 298016 70228 298072
rect 70164 298012 70228 298016
rect 71452 298012 71516 298076
rect 72556 298012 72620 298076
rect 75132 298012 75196 298076
rect 76236 298012 76300 298076
rect 77156 298072 77220 298076
rect 77156 298016 77170 298072
rect 77170 298016 77220 298072
rect 77156 298012 77220 298016
rect 78260 298012 78324 298076
rect 79732 298012 79796 298076
rect 80836 298012 80900 298076
rect 79364 297876 79428 297940
rect 80284 297876 80348 297940
rect 82124 298012 82188 298076
rect 83228 298012 83292 298076
rect 86540 298012 86604 298076
rect 87828 298012 87892 298076
rect 88932 298012 88996 298076
rect 89300 298012 89364 298076
rect 90772 298012 90836 298076
rect 93532 298012 93596 298076
rect 95004 298072 95068 298076
rect 95004 298016 95054 298072
rect 95054 298016 95068 298072
rect 95004 298012 95068 298016
rect 83044 297876 83108 297940
rect 84516 297876 84580 297940
rect 86908 297876 86972 297940
rect 87644 297876 87708 297940
rect 90220 297876 90284 297940
rect 91324 297876 91388 297940
rect 93164 297876 93228 297940
rect 94452 297876 94516 297940
rect 97028 298072 97092 298076
rect 97028 298016 97078 298072
rect 97078 298016 97092 298072
rect 97028 298012 97092 298016
rect 97948 298072 98012 298076
rect 97948 298016 97962 298072
rect 97962 298016 98012 298072
rect 97948 298012 98012 298016
rect 96660 297876 96724 297940
rect 100524 298012 100588 298076
rect 101444 298012 101508 298076
rect 104020 298012 104084 298076
rect 104388 298012 104452 298076
rect 105308 298012 105372 298076
rect 105676 298012 105740 298076
rect 106596 298072 106660 298076
rect 106596 298016 106646 298072
rect 106646 298016 106660 298072
rect 106596 298012 106660 298016
rect 106964 298012 107028 298076
rect 107700 298072 107764 298076
rect 107700 298016 107750 298072
rect 107750 298016 107764 298072
rect 107700 298012 107764 298016
rect 107884 298012 107948 298076
rect 109356 298012 109420 298076
rect 110644 298012 110708 298076
rect 113036 298072 113100 298076
rect 113036 298016 113050 298072
rect 113050 298016 113100 298072
rect 113036 298012 113100 298016
rect 114324 298012 114388 298076
rect 115612 298012 115676 298076
rect 116900 298012 116964 298076
rect 215892 298072 215956 298076
rect 215892 298016 215906 298072
rect 215906 298016 215956 298072
rect 215892 298012 215956 298016
rect 226748 298012 226812 298076
rect 227852 298012 227916 298076
rect 231348 298012 231412 298076
rect 232636 298012 232700 298076
rect 233556 298012 233620 298076
rect 235028 298012 235092 298076
rect 237236 298072 237300 298076
rect 237236 298016 237250 298072
rect 237250 298016 237300 298072
rect 237236 298012 237300 298016
rect 238340 298012 238404 298076
rect 240364 298012 240428 298076
rect 240732 298012 240796 298076
rect 242940 298072 243004 298076
rect 242940 298016 242954 298072
rect 242954 298016 243004 298072
rect 242940 298012 243004 298016
rect 244044 298072 244108 298076
rect 244044 298016 244094 298072
rect 244094 298016 244108 298072
rect 244044 298012 244108 298016
rect 244412 298012 244476 298076
rect 245516 298072 245580 298076
rect 245516 298016 245566 298072
rect 245566 298016 245580 298072
rect 245516 298012 245580 298016
rect 246804 298072 246868 298076
rect 246804 298016 246854 298072
rect 246854 298016 246868 298072
rect 246804 298012 246868 298016
rect 247908 298012 247972 298076
rect 249380 298012 249444 298076
rect 250668 298012 250732 298076
rect 252508 298012 252572 298076
rect 253612 298012 253676 298076
rect 254900 298012 254964 298076
rect 256004 298012 256068 298076
rect 259316 298012 259380 298076
rect 260788 298012 260852 298076
rect 100708 297876 100772 297940
rect 111932 297876 111996 297940
rect 237788 297876 237852 297940
rect 239260 297876 239324 297940
rect 242020 297876 242084 297940
rect 245700 297876 245764 297940
rect 247724 297876 247788 297940
rect 249012 297876 249076 297940
rect 250300 297876 250364 297940
rect 251404 297876 251468 297940
rect 253060 297876 253124 297940
rect 254532 297876 254596 297940
rect 255636 297876 255700 297940
rect 257108 297876 257172 297940
rect 259132 297876 259196 297940
rect 260604 297876 260668 297940
rect 263180 298012 263244 298076
rect 274404 298012 274468 298076
rect 276796 298012 276860 298076
rect 262996 297876 263060 297940
rect 85804 297740 85868 297804
rect 92612 297740 92676 297804
rect 101812 297740 101876 297804
rect 230060 297740 230124 297804
rect 236500 297740 236564 297804
rect 241836 297740 241900 297804
rect 246620 297740 246684 297804
rect 251956 297740 252020 297804
rect 256740 297740 256804 297804
rect 258396 297740 258460 297804
rect 99052 297468 99116 297532
rect 408540 297468 408604 297532
rect 98316 297332 98380 297396
rect 408724 297332 408788 297396
rect 83964 297060 84028 297124
rect 266860 297060 266924 297124
rect 264100 296924 264164 296988
rect 266676 296924 266740 296988
rect 264468 296788 264532 296852
rect 265756 296788 265820 296852
rect 267596 296848 267660 296852
rect 267596 296792 267610 296848
rect 267610 296792 267660 296848
rect 267596 296788 267660 296792
rect 267964 296788 268028 296852
rect 269252 296788 269316 296852
rect 270540 296788 270604 296852
rect 273116 296848 273180 296852
rect 273116 296792 273166 296848
rect 273166 296792 273180 296848
rect 273116 296788 273180 296792
rect 409276 251772 409340 251836
rect 409276 248236 409340 248300
rect 409276 237764 409340 237828
rect 409276 234228 409340 234292
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 132000 31574 140058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 132000 38414 146898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 132000 42134 150618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 381500 49574 410058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381500 56414 416898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 381500 60134 384618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 381500 63854 388338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 381500 67574 392058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 381500 74414 398898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 381500 78134 402618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 381500 81854 406338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 381500 85574 410058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381500 92414 416898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 381500 96134 384618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 381500 99854 388338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 381500 103574 392058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 381500 110414 398898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 381500 114134 402618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 381500 117854 406338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 381500 121574 410058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381500 128414 416898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 381500 132134 384618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 381500 135854 388338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 381500 139574 392058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 381500 146414 398898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 50952 363454 51300 363486
rect 50952 363218 51008 363454
rect 51244 363218 51300 363454
rect 50952 363134 51300 363218
rect 50952 362898 51008 363134
rect 51244 362898 51300 363134
rect 50952 362866 51300 362898
rect 144656 363454 145004 363486
rect 144656 363218 144712 363454
rect 144948 363218 145004 363454
rect 144656 363134 145004 363218
rect 144656 362898 144712 363134
rect 144948 362898 145004 363134
rect 144656 362866 145004 362898
rect 50272 345454 50620 345486
rect 50272 345218 50328 345454
rect 50564 345218 50620 345454
rect 50272 345134 50620 345218
rect 50272 344898 50328 345134
rect 50564 344898 50620 345134
rect 50272 344866 50620 344898
rect 145336 345454 145684 345486
rect 145336 345218 145392 345454
rect 145628 345218 145684 345454
rect 145336 345134 145684 345218
rect 145336 344898 145392 345134
rect 145628 344898 145684 345134
rect 145336 344866 145684 344898
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 50952 327454 51300 327486
rect 50952 327218 51008 327454
rect 51244 327218 51300 327454
rect 50952 327134 51300 327218
rect 50952 326898 51008 327134
rect 51244 326898 51300 327134
rect 50952 326866 51300 326898
rect 144656 327454 145004 327486
rect 144656 327218 144712 327454
rect 144948 327218 145004 327454
rect 144656 327134 145004 327218
rect 144656 326898 144712 327134
rect 144948 326898 145004 327134
rect 144656 326866 145004 326898
rect 50272 309454 50620 309486
rect 50272 309218 50328 309454
rect 50564 309218 50620 309454
rect 50272 309134 50620 309218
rect 50272 308898 50328 309134
rect 50564 308898 50620 309134
rect 50272 308866 50620 308898
rect 145336 309454 145684 309486
rect 145336 309218 145392 309454
rect 145628 309218 145684 309454
rect 145336 309134 145684 309218
rect 145336 308898 145392 309134
rect 145628 308898 145684 309134
rect 145336 308866 145684 308898
rect 55856 299573 55916 300106
rect 55853 299572 55919 299573
rect 55853 299508 55854 299572
rect 55918 299508 55919 299572
rect 65512 299570 65572 300106
rect 66736 299570 66796 300106
rect 67824 299573 67884 300106
rect 65512 299510 65626 299570
rect 55853 299507 55919 299508
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 65566 298077 65626 299510
rect 66670 299510 66796 299570
rect 67821 299572 67887 299573
rect 66670 298077 66730 299510
rect 67821 299508 67822 299572
rect 67886 299508 67887 299572
rect 69184 299570 69244 300106
rect 70136 299570 70196 300106
rect 71360 299570 71420 300106
rect 72584 299570 72644 300106
rect 73672 299570 73732 300106
rect 69184 299510 69306 299570
rect 70136 299510 70226 299570
rect 71360 299510 71514 299570
rect 67821 299507 67887 299508
rect 69246 298077 69306 299510
rect 70166 298077 70226 299510
rect 71454 298077 71514 299510
rect 72558 299510 72644 299570
rect 73662 299510 73732 299570
rect 75032 299570 75092 300106
rect 76120 299570 76180 300106
rect 77208 299570 77268 300106
rect 75032 299510 75194 299570
rect 76120 299510 76298 299570
rect 72558 298077 72618 299510
rect 73662 298213 73722 299510
rect 73659 298212 73725 298213
rect 73659 298148 73660 298212
rect 73724 298148 73725 298212
rect 73659 298147 73725 298148
rect 75134 298077 75194 299510
rect 76238 298077 76298 299510
rect 77158 299510 77268 299570
rect 77888 299570 77948 300106
rect 78296 299570 78356 300106
rect 77888 299510 77954 299570
rect 77158 298077 77218 299510
rect 77894 298213 77954 299510
rect 78262 299510 78356 299570
rect 79248 299570 79308 300106
rect 79656 299570 79716 300106
rect 80336 299570 80396 300106
rect 79248 299510 79426 299570
rect 79656 299510 79794 299570
rect 77891 298212 77957 298213
rect 77891 298148 77892 298212
rect 77956 298148 77957 298212
rect 77891 298147 77957 298148
rect 78262 298077 78322 299510
rect 65563 298076 65629 298077
rect 65563 298012 65564 298076
rect 65628 298012 65629 298076
rect 65563 298011 65629 298012
rect 66667 298076 66733 298077
rect 66667 298012 66668 298076
rect 66732 298012 66733 298076
rect 66667 298011 66733 298012
rect 69243 298076 69309 298077
rect 69243 298012 69244 298076
rect 69308 298012 69309 298076
rect 69243 298011 69309 298012
rect 70163 298076 70229 298077
rect 70163 298012 70164 298076
rect 70228 298012 70229 298076
rect 70163 298011 70229 298012
rect 71451 298076 71517 298077
rect 71451 298012 71452 298076
rect 71516 298012 71517 298076
rect 71451 298011 71517 298012
rect 72555 298076 72621 298077
rect 72555 298012 72556 298076
rect 72620 298012 72621 298076
rect 72555 298011 72621 298012
rect 75131 298076 75197 298077
rect 75131 298012 75132 298076
rect 75196 298012 75197 298076
rect 75131 298011 75197 298012
rect 76235 298076 76301 298077
rect 76235 298012 76236 298076
rect 76300 298012 76301 298076
rect 76235 298011 76301 298012
rect 77155 298076 77221 298077
rect 77155 298012 77156 298076
rect 77220 298012 77221 298076
rect 77155 298011 77221 298012
rect 78259 298076 78325 298077
rect 78259 298012 78260 298076
rect 78324 298012 78325 298076
rect 78259 298011 78325 298012
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 132000 45854 154338
rect 48954 266614 49574 298000
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 132000 49574 158058
rect 55794 273454 56414 298000
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 132000 56414 164898
rect 59514 277174 60134 298000
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 132000 60134 132618
rect 63234 280894 63854 298000
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 132000 63854 136338
rect 66954 284614 67574 298000
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 132000 67574 140058
rect 73794 291454 74414 298000
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 132000 74414 146898
rect 77514 295174 78134 298000
rect 79366 297941 79426 299510
rect 79734 298077 79794 299510
rect 80286 299510 80396 299570
rect 80744 299570 80804 300106
rect 81832 299570 81892 300106
rect 80744 299510 80898 299570
rect 79731 298076 79797 298077
rect 79731 298012 79732 298076
rect 79796 298012 79797 298076
rect 79731 298011 79797 298012
rect 80286 297941 80346 299510
rect 80838 298077 80898 299510
rect 81758 299510 81892 299570
rect 81968 299570 82028 300106
rect 83056 299570 83116 300106
rect 81968 299510 82186 299570
rect 81758 298213 81818 299510
rect 81755 298212 81821 298213
rect 81755 298148 81756 298212
rect 81820 298148 81821 298212
rect 81755 298147 81821 298148
rect 82126 298077 82186 299510
rect 83046 299510 83116 299570
rect 83192 299570 83252 300106
rect 84144 299570 84204 300106
rect 83192 299510 83290 299570
rect 80835 298076 80901 298077
rect 80835 298012 80836 298076
rect 80900 298012 80901 298076
rect 80835 298011 80901 298012
rect 82123 298076 82189 298077
rect 82123 298012 82124 298076
rect 82188 298012 82189 298076
rect 82123 298011 82189 298012
rect 79363 297940 79429 297941
rect 79363 297876 79364 297940
rect 79428 297876 79429 297940
rect 79363 297875 79429 297876
rect 80283 297940 80349 297941
rect 80283 297876 80284 297940
rect 80348 297876 80349 297940
rect 80283 297875 80349 297876
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 132000 78134 150618
rect 81234 262894 81854 298000
rect 83046 297941 83106 299510
rect 83230 298077 83290 299510
rect 83966 299510 84204 299570
rect 84416 299570 84476 300106
rect 85504 299570 85564 300106
rect 84416 299510 84578 299570
rect 83227 298076 83293 298077
rect 83227 298012 83228 298076
rect 83292 298012 83293 298076
rect 83227 298011 83293 298012
rect 83043 297940 83109 297941
rect 83043 297876 83044 297940
rect 83108 297876 83109 297940
rect 83043 297875 83109 297876
rect 83966 297125 84026 299510
rect 84518 297941 84578 299510
rect 85438 299510 85564 299570
rect 85640 299570 85700 300106
rect 86592 299570 86652 300106
rect 85640 299510 85866 299570
rect 85438 298213 85498 299510
rect 85435 298212 85501 298213
rect 85435 298148 85436 298212
rect 85500 298148 85501 298212
rect 85435 298147 85501 298148
rect 84515 297940 84581 297941
rect 84515 297876 84516 297940
rect 84580 297876 84581 297940
rect 84515 297875 84581 297876
rect 83963 297124 84029 297125
rect 83963 297060 83964 297124
rect 84028 297060 84029 297124
rect 83963 297059 84029 297060
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 132000 81854 154338
rect 84954 266614 85574 298000
rect 85806 297805 85866 299510
rect 86542 299510 86652 299570
rect 86864 299570 86924 300106
rect 87680 299570 87740 300106
rect 86864 299510 86970 299570
rect 86542 298077 86602 299510
rect 86539 298076 86605 298077
rect 86539 298012 86540 298076
rect 86604 298012 86605 298076
rect 86539 298011 86605 298012
rect 86910 297941 86970 299510
rect 87646 299510 87740 299570
rect 87816 299570 87876 300106
rect 88904 299570 88964 300106
rect 89312 299570 89372 300106
rect 90264 299570 90324 300106
rect 87816 299510 87890 299570
rect 88904 299510 88994 299570
rect 87646 297941 87706 299510
rect 87830 298077 87890 299510
rect 88934 298077 88994 299510
rect 89302 299510 89372 299570
rect 90222 299510 90324 299570
rect 90672 299570 90732 300106
rect 91352 299570 91412 300106
rect 91896 299570 91956 300106
rect 90672 299510 90834 299570
rect 89302 298077 89362 299510
rect 87827 298076 87893 298077
rect 87827 298012 87828 298076
rect 87892 298012 87893 298076
rect 87827 298011 87893 298012
rect 88931 298076 88997 298077
rect 88931 298012 88932 298076
rect 88996 298012 88997 298076
rect 88931 298011 88997 298012
rect 89299 298076 89365 298077
rect 89299 298012 89300 298076
rect 89364 298012 89365 298076
rect 89299 298011 89365 298012
rect 90222 297941 90282 299510
rect 90774 298077 90834 299510
rect 91326 299510 91412 299570
rect 91878 299510 91956 299570
rect 92440 299570 92500 300106
rect 93120 299570 93180 300106
rect 93528 299570 93588 300106
rect 94344 299842 94404 300106
rect 94888 299842 94948 300106
rect 94344 299782 94514 299842
rect 94888 299782 95066 299842
rect 92440 299510 92674 299570
rect 93120 299510 93226 299570
rect 93528 299510 93594 299570
rect 90771 298076 90837 298077
rect 90771 298012 90772 298076
rect 90836 298012 90837 298076
rect 90771 298011 90837 298012
rect 91326 297941 91386 299510
rect 91878 298213 91938 299510
rect 91875 298212 91941 298213
rect 91875 298148 91876 298212
rect 91940 298148 91941 298212
rect 91875 298147 91941 298148
rect 86907 297940 86973 297941
rect 86907 297876 86908 297940
rect 86972 297876 86973 297940
rect 86907 297875 86973 297876
rect 87643 297940 87709 297941
rect 87643 297876 87644 297940
rect 87708 297876 87709 297940
rect 87643 297875 87709 297876
rect 90219 297940 90285 297941
rect 90219 297876 90220 297940
rect 90284 297876 90285 297940
rect 90219 297875 90285 297876
rect 91323 297940 91389 297941
rect 91323 297876 91324 297940
rect 91388 297876 91389 297940
rect 91323 297875 91389 297876
rect 85803 297804 85869 297805
rect 85803 297740 85804 297804
rect 85868 297740 85869 297804
rect 85803 297739 85869 297740
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 132000 85574 158058
rect 91794 273454 92414 298000
rect 92614 297805 92674 299510
rect 93166 297941 93226 299510
rect 93534 298077 93594 299510
rect 93531 298076 93597 298077
rect 93531 298012 93532 298076
rect 93596 298012 93597 298076
rect 93531 298011 93597 298012
rect 94454 297941 94514 299782
rect 95006 298077 95066 299782
rect 95568 299570 95628 300106
rect 95976 299570 96036 300106
rect 95558 299510 95628 299570
rect 95926 299510 96036 299570
rect 96656 299570 96716 300106
rect 97064 299570 97124 300106
rect 97880 299842 97940 300106
rect 97880 299782 98010 299842
rect 96656 299510 96722 299570
rect 95558 298213 95618 299510
rect 95926 298213 95986 299510
rect 95555 298212 95621 298213
rect 95555 298148 95556 298212
rect 95620 298148 95621 298212
rect 95555 298147 95621 298148
rect 95923 298212 95989 298213
rect 95923 298148 95924 298212
rect 95988 298148 95989 298212
rect 95923 298147 95989 298148
rect 95003 298076 95069 298077
rect 95003 298012 95004 298076
rect 95068 298012 95069 298076
rect 95003 298011 95069 298012
rect 93163 297940 93229 297941
rect 93163 297876 93164 297940
rect 93228 297876 93229 297940
rect 93163 297875 93229 297876
rect 94451 297940 94517 297941
rect 94451 297876 94452 297940
rect 94516 297876 94517 297940
rect 94451 297875 94517 297876
rect 92611 297804 92677 297805
rect 92611 297740 92612 297804
rect 92676 297740 92677 297804
rect 92611 297739 92677 297740
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 132000 92414 164898
rect 95514 277174 96134 298000
rect 96662 297941 96722 299510
rect 97030 299510 97124 299570
rect 97030 298077 97090 299510
rect 97950 298077 98010 299782
rect 98288 299570 98348 300106
rect 99104 299570 99164 300106
rect 98288 299510 98378 299570
rect 97027 298076 97093 298077
rect 97027 298012 97028 298076
rect 97092 298012 97093 298076
rect 97027 298011 97093 298012
rect 97947 298076 98013 298077
rect 97947 298012 97948 298076
rect 98012 298012 98013 298076
rect 97947 298011 98013 298012
rect 96659 297940 96725 297941
rect 96659 297876 96660 297940
rect 96724 297876 96725 297940
rect 96659 297875 96725 297876
rect 98318 297397 98378 299510
rect 99054 299510 99164 299570
rect 99376 299570 99436 300106
rect 100600 299842 100660 300106
rect 100526 299782 100660 299842
rect 99376 299510 99482 299570
rect 99054 297533 99114 299510
rect 99422 298213 99482 299510
rect 99419 298212 99485 298213
rect 99419 298148 99420 298212
rect 99484 298148 99485 298212
rect 99419 298147 99485 298148
rect 100526 298077 100586 299782
rect 100736 299570 100796 300106
rect 100710 299510 100796 299570
rect 101416 299570 101476 300106
rect 101824 299570 101884 300106
rect 101416 299510 101506 299570
rect 100523 298076 100589 298077
rect 100523 298012 100524 298076
rect 100588 298012 100589 298076
rect 100523 298011 100589 298012
rect 99051 297532 99117 297533
rect 99051 297468 99052 297532
rect 99116 297468 99117 297532
rect 99051 297467 99117 297468
rect 98315 297396 98381 297397
rect 98315 297332 98316 297396
rect 98380 297332 98381 297396
rect 98315 297331 98381 297332
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 132000 96134 132618
rect 99234 280894 99854 298000
rect 100710 297941 100770 299510
rect 101446 298077 101506 299510
rect 101814 299510 101884 299570
rect 102912 299570 102972 300106
rect 103184 299842 103244 300106
rect 103184 299782 103346 299842
rect 102912 299510 102978 299570
rect 101443 298076 101509 298077
rect 101443 298012 101444 298076
rect 101508 298012 101509 298076
rect 101443 298011 101509 298012
rect 100707 297940 100773 297941
rect 100707 297876 100708 297940
rect 100772 297876 100773 297940
rect 100707 297875 100773 297876
rect 101814 297805 101874 299510
rect 102918 298213 102978 299510
rect 103286 298213 103346 299782
rect 104000 299570 104060 300106
rect 104408 299570 104468 300106
rect 105224 299842 105284 300106
rect 105224 299782 105370 299842
rect 104000 299510 104082 299570
rect 102915 298212 102981 298213
rect 102915 298148 102916 298212
rect 102980 298148 102981 298212
rect 102915 298147 102981 298148
rect 103283 298212 103349 298213
rect 103283 298148 103284 298212
rect 103348 298148 103349 298212
rect 103283 298147 103349 298148
rect 104022 298077 104082 299510
rect 104390 299510 104468 299570
rect 104390 298077 104450 299510
rect 105310 298077 105370 299782
rect 105632 299570 105692 300106
rect 106584 299570 106644 300106
rect 106856 299842 106916 300106
rect 106856 299782 107026 299842
rect 105632 299510 105738 299570
rect 106584 299510 106658 299570
rect 105678 298077 105738 299510
rect 106598 298077 106658 299510
rect 106966 298077 107026 299782
rect 107672 299570 107732 300106
rect 107808 299842 107868 300106
rect 107808 299782 107946 299842
rect 107672 299510 107762 299570
rect 107702 298077 107762 299510
rect 107886 298077 107946 299782
rect 109304 299570 109364 300106
rect 110528 299842 110588 300106
rect 110528 299782 110706 299842
rect 109304 299510 109418 299570
rect 109358 298077 109418 299510
rect 110646 298077 110706 299782
rect 111888 299570 111948 300106
rect 113112 299842 113172 300106
rect 113038 299782 113172 299842
rect 111888 299510 111994 299570
rect 104019 298076 104085 298077
rect 104019 298012 104020 298076
rect 104084 298012 104085 298076
rect 104019 298011 104085 298012
rect 104387 298076 104453 298077
rect 104387 298012 104388 298076
rect 104452 298012 104453 298076
rect 104387 298011 104453 298012
rect 105307 298076 105373 298077
rect 105307 298012 105308 298076
rect 105372 298012 105373 298076
rect 105307 298011 105373 298012
rect 105675 298076 105741 298077
rect 105675 298012 105676 298076
rect 105740 298012 105741 298076
rect 105675 298011 105741 298012
rect 106595 298076 106661 298077
rect 106595 298012 106596 298076
rect 106660 298012 106661 298076
rect 106595 298011 106661 298012
rect 106963 298076 107029 298077
rect 106963 298012 106964 298076
rect 107028 298012 107029 298076
rect 106963 298011 107029 298012
rect 107699 298076 107765 298077
rect 107699 298012 107700 298076
rect 107764 298012 107765 298076
rect 107699 298011 107765 298012
rect 107883 298076 107949 298077
rect 107883 298012 107884 298076
rect 107948 298012 107949 298076
rect 107883 298011 107949 298012
rect 109355 298076 109421 298077
rect 109355 298012 109356 298076
rect 109420 298012 109421 298076
rect 109355 298011 109421 298012
rect 110643 298076 110709 298077
rect 110643 298012 110644 298076
rect 110708 298012 110709 298076
rect 110643 298011 110709 298012
rect 101811 297804 101877 297805
rect 101811 297740 101812 297804
rect 101876 297740 101877 297804
rect 101811 297739 101877 297740
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 132000 99854 136338
rect 102954 284614 103574 298000
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 132000 103574 140058
rect 109794 291454 110414 298000
rect 111934 297941 111994 299510
rect 113038 298077 113098 299782
rect 114336 299570 114396 300106
rect 114326 299510 114396 299570
rect 115560 299570 115620 300106
rect 116784 299570 116844 300106
rect 115560 299510 115674 299570
rect 116784 299510 116962 299570
rect 114326 298077 114386 299510
rect 115614 298077 115674 299510
rect 116902 298077 116962 299510
rect 113035 298076 113101 298077
rect 113035 298012 113036 298076
rect 113100 298012 113101 298076
rect 113035 298011 113101 298012
rect 114323 298076 114389 298077
rect 114323 298012 114324 298076
rect 114388 298012 114389 298076
rect 114323 298011 114389 298012
rect 115611 298076 115677 298077
rect 115611 298012 115612 298076
rect 115676 298012 115677 298076
rect 115611 298011 115677 298012
rect 116899 298076 116965 298077
rect 116899 298012 116900 298076
rect 116964 298012 116965 298076
rect 116899 298011 116965 298012
rect 111931 297940 111997 297941
rect 111931 297876 111932 297940
rect 111996 297876 111997 297940
rect 111931 297875 111997 297876
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 132000 110414 146898
rect 113514 295174 114134 298000
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 132000 114134 150618
rect 117234 262894 117854 298000
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 132000 117854 154338
rect 120954 266614 121574 298000
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 132000 121574 158058
rect 127794 273454 128414 298000
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 132000 128414 164898
rect 131514 277174 132134 298000
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 132000 132134 132618
rect 135234 280894 135854 298000
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 34208 111454 34528 111486
rect 34208 111218 34250 111454
rect 34486 111218 34528 111454
rect 34208 111134 34528 111218
rect 34208 110898 34250 111134
rect 34486 110898 34528 111134
rect 34208 110866 34528 110898
rect 64928 111454 65248 111486
rect 64928 111218 64970 111454
rect 65206 111218 65248 111454
rect 64928 111134 65248 111218
rect 64928 110898 64970 111134
rect 65206 110898 65248 111134
rect 64928 110866 65248 110898
rect 95648 111454 95968 111486
rect 95648 111218 95690 111454
rect 95926 111218 95968 111454
rect 95648 111134 95968 111218
rect 95648 110898 95690 111134
rect 95926 110898 95968 111134
rect 95648 110866 95968 110898
rect 126368 111454 126688 111486
rect 126368 111218 126410 111454
rect 126646 111218 126688 111454
rect 126368 111134 126688 111218
rect 126368 110898 126410 111134
rect 126646 110898 126688 111134
rect 126368 110866 126688 110898
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 49568 93454 49888 93486
rect 49568 93218 49610 93454
rect 49846 93218 49888 93454
rect 49568 93134 49888 93218
rect 49568 92898 49610 93134
rect 49846 92898 49888 93134
rect 49568 92866 49888 92898
rect 80288 93454 80608 93486
rect 80288 93218 80330 93454
rect 80566 93218 80608 93454
rect 80288 93134 80608 93218
rect 80288 92898 80330 93134
rect 80566 92898 80608 93134
rect 80288 92866 80608 92898
rect 111008 93454 111328 93486
rect 111008 93218 111050 93454
rect 111286 93218 111328 93454
rect 111008 93134 111328 93218
rect 111008 92898 111050 93134
rect 111286 92898 111328 93134
rect 111008 92866 111328 92898
rect 34208 75454 34528 75486
rect 34208 75218 34250 75454
rect 34486 75218 34528 75454
rect 34208 75134 34528 75218
rect 34208 74898 34250 75134
rect 34486 74898 34528 75134
rect 34208 74866 34528 74898
rect 64928 75454 65248 75486
rect 64928 75218 64970 75454
rect 65206 75218 65248 75454
rect 64928 75134 65248 75218
rect 64928 74898 64970 75134
rect 65206 74898 65248 75134
rect 64928 74866 65248 74898
rect 95648 75454 95968 75486
rect 95648 75218 95690 75454
rect 95926 75218 95968 75454
rect 95648 75134 95968 75218
rect 95648 74898 95690 75134
rect 95926 74898 95968 75134
rect 95648 74866 95968 74898
rect 126368 75454 126688 75486
rect 126368 75218 126410 75454
rect 126646 75218 126688 75454
rect 126368 75134 126688 75218
rect 126368 74898 126410 75134
rect 126646 74898 126688 75134
rect 126368 74866 126688 74898
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 49568 57454 49888 57486
rect 49568 57218 49610 57454
rect 49846 57218 49888 57454
rect 49568 57134 49888 57218
rect 49568 56898 49610 57134
rect 49846 56898 49888 57134
rect 49568 56866 49888 56898
rect 80288 57454 80608 57486
rect 80288 57218 80330 57454
rect 80566 57218 80608 57454
rect 80288 57134 80608 57218
rect 80288 56898 80330 57134
rect 80566 56898 80608 57134
rect 80288 56866 80608 56898
rect 111008 57454 111328 57486
rect 111008 57218 111050 57454
rect 111286 57218 111328 57454
rect 111008 57134 111328 57218
rect 111008 56898 111050 57134
rect 111286 56898 111328 57134
rect 111008 56866 111328 56898
rect 34208 39454 34528 39486
rect 34208 39218 34250 39454
rect 34486 39218 34528 39454
rect 34208 39134 34528 39218
rect 34208 38898 34250 39134
rect 34486 38898 34528 39134
rect 34208 38866 34528 38898
rect 64928 39454 65248 39486
rect 64928 39218 64970 39454
rect 65206 39218 65248 39454
rect 64928 39134 65248 39218
rect 64928 38898 64970 39134
rect 65206 38898 65248 39134
rect 64928 38866 65248 38898
rect 95648 39454 95968 39486
rect 95648 39218 95690 39454
rect 95926 39218 95968 39454
rect 95648 39134 95968 39218
rect 95648 38898 95690 39134
rect 95926 38898 95968 39134
rect 95648 38866 95968 38898
rect 126368 39454 126688 39486
rect 126368 39218 126410 39454
rect 126646 39218 126688 39454
rect 126368 39134 126688 39218
rect 126368 38898 126410 39134
rect 126646 38898 126688 39134
rect 126368 38866 126688 38898
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 28000
rect 37794 3454 38414 28000
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 7174 42134 28000
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 10894 45854 28000
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 14614 49574 28000
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 28000
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 28000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 28000
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 28000
rect 73794 3454 74414 28000
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 7174 78134 28000
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 10894 81854 28000
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 14614 85574 28000
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 21454 92414 28000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 28000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 -5146 99854 28000
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 28000
rect 109794 3454 110414 28000
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 7174 114134 28000
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 10894 117854 28000
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 14614 121574 28000
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 21454 128414 28000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 28000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 284614 139574 298000
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 291454 146414 298000
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 252000 189854 262338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 252000 193574 266058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 252000 200414 272898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 252000 204134 276618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 381500 211574 392058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 381500 218414 398898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 381500 222134 402618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 381500 225854 406338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 381500 229574 410058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381500 236414 416898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 381500 240134 384618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 381500 243854 388338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 381500 247574 392058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 381500 254414 398898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 381500 258134 402618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 381500 261854 406338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 381500 265574 410058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381500 272414 416898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 381500 276134 384618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 381500 279854 388338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 381500 283574 392058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 381500 290414 398898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 381500 294134 402618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 381500 297854 406338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 381500 301574 410058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381500 308414 416898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 210952 363454 211300 363486
rect 210952 363218 211008 363454
rect 211244 363218 211300 363454
rect 210952 363134 211300 363218
rect 210952 362898 211008 363134
rect 211244 362898 211300 363134
rect 210952 362866 211300 362898
rect 304656 363454 305004 363486
rect 304656 363218 304712 363454
rect 304948 363218 305004 363454
rect 304656 363134 305004 363218
rect 304656 362898 304712 363134
rect 304948 362898 305004 363134
rect 304656 362866 305004 362898
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 210272 345454 210620 345486
rect 210272 345218 210328 345454
rect 210564 345218 210620 345454
rect 210272 345134 210620 345218
rect 210272 344898 210328 345134
rect 210564 344898 210620 345134
rect 210272 344866 210620 344898
rect 305336 345454 305684 345486
rect 305336 345218 305392 345454
rect 305628 345218 305684 345454
rect 305336 345134 305684 345218
rect 305336 344898 305392 345134
rect 305628 344898 305684 345134
rect 305336 344866 305684 344898
rect 210952 327454 211300 327486
rect 210952 327218 211008 327454
rect 211244 327218 211300 327454
rect 210952 327134 211300 327218
rect 210952 326898 211008 327134
rect 211244 326898 211300 327134
rect 210952 326866 211300 326898
rect 304656 327454 305004 327486
rect 304656 327218 304712 327454
rect 304948 327218 305004 327454
rect 304656 327134 305004 327218
rect 304656 326898 304712 327134
rect 304948 326898 305004 327134
rect 304656 326866 305004 326898
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 210272 309454 210620 309486
rect 210272 309218 210328 309454
rect 210564 309218 210620 309454
rect 210272 309134 210620 309218
rect 210272 308898 210328 309134
rect 210564 308898 210620 309134
rect 210272 308866 210620 308898
rect 305336 309454 305684 309486
rect 305336 309218 305392 309454
rect 305628 309218 305684 309454
rect 305336 309134 305684 309218
rect 305336 308898 305392 309134
rect 305628 308898 305684 309134
rect 305336 308866 305684 308898
rect 215856 299570 215916 300106
rect 225512 299570 225572 300106
rect 215856 299510 215954 299570
rect 215894 298077 215954 299510
rect 225462 299510 225572 299570
rect 226736 299570 226796 300106
rect 227824 299570 227884 300106
rect 229184 299570 229244 300106
rect 230136 299570 230196 300106
rect 231360 299570 231420 300106
rect 226736 299510 226810 299570
rect 227824 299510 227914 299570
rect 225462 298213 225522 299510
rect 225459 298212 225525 298213
rect 225459 298148 225460 298212
rect 225524 298148 225525 298212
rect 225459 298147 225525 298148
rect 226750 298077 226810 299510
rect 227854 298077 227914 299510
rect 229142 299510 229244 299570
rect 230062 299510 230196 299570
rect 231350 299510 231420 299570
rect 232584 299570 232644 300106
rect 233672 299570 233732 300106
rect 235032 299570 235092 300106
rect 232584 299510 232698 299570
rect 229142 298349 229202 299510
rect 229139 298348 229205 298349
rect 229139 298284 229140 298348
rect 229204 298284 229205 298348
rect 229139 298283 229205 298284
rect 215891 298076 215957 298077
rect 215891 298012 215892 298076
rect 215956 298012 215957 298076
rect 215891 298011 215957 298012
rect 226747 298076 226813 298077
rect 226747 298012 226748 298076
rect 226812 298012 226813 298076
rect 226747 298011 226813 298012
rect 227851 298076 227917 298077
rect 227851 298012 227852 298076
rect 227916 298012 227917 298076
rect 227851 298011 227917 298012
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 252000 207854 280338
rect 210954 284614 211574 298000
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 252000 211574 284058
rect 217794 291454 218414 298000
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 252000 218414 254898
rect 221514 295174 222134 298000
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 252000 222134 258618
rect 225234 262894 225854 298000
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 252000 225854 262338
rect 228954 266614 229574 298000
rect 230062 297805 230122 299510
rect 231350 298077 231410 299510
rect 232638 298077 232698 299510
rect 233558 299510 233732 299570
rect 235030 299510 235092 299570
rect 236120 299570 236180 300106
rect 237208 299570 237268 300106
rect 237888 299570 237948 300106
rect 236120 299510 236562 299570
rect 237208 299510 237298 299570
rect 233558 298077 233618 299510
rect 235030 298077 235090 299510
rect 231347 298076 231413 298077
rect 231347 298012 231348 298076
rect 231412 298012 231413 298076
rect 231347 298011 231413 298012
rect 232635 298076 232701 298077
rect 232635 298012 232636 298076
rect 232700 298012 232701 298076
rect 232635 298011 232701 298012
rect 233555 298076 233621 298077
rect 233555 298012 233556 298076
rect 233620 298012 233621 298076
rect 233555 298011 233621 298012
rect 235027 298076 235093 298077
rect 235027 298012 235028 298076
rect 235092 298012 235093 298076
rect 235027 298011 235093 298012
rect 230059 297804 230125 297805
rect 230059 297740 230060 297804
rect 230124 297740 230125 297804
rect 230059 297739 230125 297740
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 252000 229574 266058
rect 235794 273454 236414 298000
rect 236502 297805 236562 299510
rect 237238 298077 237298 299510
rect 237790 299510 237948 299570
rect 238296 299570 238356 300106
rect 239248 299570 239308 300106
rect 239656 299845 239716 300106
rect 239653 299844 239719 299845
rect 239653 299780 239654 299844
rect 239718 299780 239719 299844
rect 239653 299779 239719 299780
rect 240336 299570 240396 300106
rect 240744 299570 240804 300106
rect 238296 299510 238402 299570
rect 239248 299510 239322 299570
rect 240336 299510 240426 299570
rect 237235 298076 237301 298077
rect 237235 298012 237236 298076
rect 237300 298012 237301 298076
rect 237235 298011 237301 298012
rect 237790 297941 237850 299510
rect 238342 298077 238402 299510
rect 238339 298076 238405 298077
rect 238339 298012 238340 298076
rect 238404 298012 238405 298076
rect 238339 298011 238405 298012
rect 239262 297941 239322 299510
rect 240366 298077 240426 299510
rect 240734 299510 240804 299570
rect 241832 299570 241892 300106
rect 241968 299570 242028 300106
rect 243056 299709 243116 300106
rect 243053 299708 243119 299709
rect 243053 299644 243054 299708
rect 243118 299644 243119 299708
rect 243053 299643 243119 299644
rect 243192 299570 243252 300106
rect 244144 299570 244204 300106
rect 244416 299570 244476 300106
rect 241832 299510 241898 299570
rect 241968 299510 242082 299570
rect 240734 298077 240794 299510
rect 240363 298076 240429 298077
rect 240363 298012 240364 298076
rect 240428 298012 240429 298076
rect 240363 298011 240429 298012
rect 240731 298076 240797 298077
rect 240731 298012 240732 298076
rect 240796 298012 240797 298076
rect 240731 298011 240797 298012
rect 237787 297940 237853 297941
rect 237787 297876 237788 297940
rect 237852 297876 237853 297940
rect 237787 297875 237853 297876
rect 239259 297940 239325 297941
rect 239259 297876 239260 297940
rect 239324 297876 239325 297940
rect 239259 297875 239325 297876
rect 236499 297804 236565 297805
rect 236499 297740 236500 297804
rect 236564 297740 236565 297804
rect 236499 297739 236565 297740
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 252000 236414 272898
rect 239514 277174 240134 298000
rect 241838 297805 241898 299510
rect 242022 297941 242082 299510
rect 242942 299510 243252 299570
rect 244046 299510 244204 299570
rect 244414 299510 244476 299570
rect 245504 299570 245564 300106
rect 245640 299570 245700 300106
rect 246592 299570 246652 300106
rect 246864 299570 246924 300106
rect 247680 299570 247740 300106
rect 245504 299510 245578 299570
rect 245640 299510 245762 299570
rect 246592 299510 246682 299570
rect 242942 298077 243002 299510
rect 244046 298077 244106 299510
rect 244414 298077 244474 299510
rect 245518 298077 245578 299510
rect 242939 298076 243005 298077
rect 242939 298012 242940 298076
rect 243004 298012 243005 298076
rect 242939 298011 243005 298012
rect 244043 298076 244109 298077
rect 244043 298012 244044 298076
rect 244108 298012 244109 298076
rect 244043 298011 244109 298012
rect 244411 298076 244477 298077
rect 244411 298012 244412 298076
rect 244476 298012 244477 298076
rect 244411 298011 244477 298012
rect 245515 298076 245581 298077
rect 245515 298012 245516 298076
rect 245580 298012 245581 298076
rect 245515 298011 245581 298012
rect 242019 297940 242085 297941
rect 242019 297876 242020 297940
rect 242084 297876 242085 297940
rect 242019 297875 242085 297876
rect 241835 297804 241901 297805
rect 241835 297740 241836 297804
rect 241900 297740 241901 297804
rect 241835 297739 241901 297740
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 252000 240134 276618
rect 243234 280894 243854 298000
rect 245702 297941 245762 299510
rect 245699 297940 245765 297941
rect 245699 297876 245700 297940
rect 245764 297876 245765 297940
rect 245699 297875 245765 297876
rect 246622 297805 246682 299510
rect 246806 299510 246924 299570
rect 247542 299510 247740 299570
rect 247816 299570 247876 300106
rect 248904 299842 248964 300106
rect 249312 299842 249372 300106
rect 248904 299782 249074 299842
rect 249312 299782 249442 299842
rect 247816 299510 247970 299570
rect 246806 298077 246866 299510
rect 247542 298890 247602 299510
rect 247542 298830 247786 298890
rect 246803 298076 246869 298077
rect 246803 298012 246804 298076
rect 246868 298012 246869 298076
rect 246803 298011 246869 298012
rect 246619 297804 246685 297805
rect 246619 297740 246620 297804
rect 246684 297740 246685 297804
rect 246619 297739 246685 297740
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 252000 243854 280338
rect 246954 284614 247574 298000
rect 247726 297941 247786 298830
rect 247910 298077 247970 299510
rect 247907 298076 247973 298077
rect 247907 298012 247908 298076
rect 247972 298012 247973 298076
rect 247907 298011 247973 298012
rect 249014 297941 249074 299782
rect 249382 298077 249442 299782
rect 250264 299570 250324 300106
rect 250672 299570 250732 300106
rect 250264 299510 250362 299570
rect 249379 298076 249445 298077
rect 249379 298012 249380 298076
rect 249444 298012 249445 298076
rect 249379 298011 249445 298012
rect 250302 297941 250362 299510
rect 250670 299510 250732 299570
rect 251352 299570 251412 300106
rect 251896 299570 251956 300106
rect 252440 299842 252500 300106
rect 252440 299782 252570 299842
rect 251352 299510 251466 299570
rect 251896 299510 252018 299570
rect 250670 298077 250730 299510
rect 250667 298076 250733 298077
rect 250667 298012 250668 298076
rect 250732 298012 250733 298076
rect 250667 298011 250733 298012
rect 251406 297941 251466 299510
rect 247723 297940 247789 297941
rect 247723 297876 247724 297940
rect 247788 297876 247789 297940
rect 247723 297875 247789 297876
rect 249011 297940 249077 297941
rect 249011 297876 249012 297940
rect 249076 297876 249077 297940
rect 249011 297875 249077 297876
rect 250299 297940 250365 297941
rect 250299 297876 250300 297940
rect 250364 297876 250365 297940
rect 250299 297875 250365 297876
rect 251403 297940 251469 297941
rect 251403 297876 251404 297940
rect 251468 297876 251469 297940
rect 251403 297875 251469 297876
rect 251958 297805 252018 299510
rect 252510 298077 252570 299782
rect 253120 299570 253180 300106
rect 253528 299842 253588 300106
rect 253528 299782 253674 299842
rect 253062 299510 253180 299570
rect 252507 298076 252573 298077
rect 252507 298012 252508 298076
rect 252572 298012 252573 298076
rect 252507 298011 252573 298012
rect 253062 297941 253122 299510
rect 253614 298077 253674 299782
rect 254344 299570 254404 300106
rect 254888 299570 254948 300106
rect 255568 299842 255628 300106
rect 255568 299782 255698 299842
rect 254344 299510 254594 299570
rect 254888 299510 254962 299570
rect 253611 298076 253677 298077
rect 253611 298012 253612 298076
rect 253676 298012 253677 298076
rect 253611 298011 253677 298012
rect 253059 297940 253125 297941
rect 253059 297876 253060 297940
rect 253124 297876 253125 297940
rect 253059 297875 253125 297876
rect 251955 297804 252021 297805
rect 251955 297740 251956 297804
rect 252020 297740 252021 297804
rect 251955 297739 252021 297740
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 252000 247574 284058
rect 253794 291454 254414 298000
rect 254534 297941 254594 299510
rect 254902 298077 254962 299510
rect 254899 298076 254965 298077
rect 254899 298012 254900 298076
rect 254964 298012 254965 298076
rect 254899 298011 254965 298012
rect 255638 297941 255698 299782
rect 255976 299570 256036 300106
rect 256656 299842 256716 300106
rect 256656 299782 256802 299842
rect 255976 299510 256066 299570
rect 256006 298077 256066 299510
rect 256003 298076 256069 298077
rect 256003 298012 256004 298076
rect 256068 298012 256069 298076
rect 256003 298011 256069 298012
rect 254531 297940 254597 297941
rect 254531 297876 254532 297940
rect 254596 297876 254597 297940
rect 254531 297875 254597 297876
rect 255635 297940 255701 297941
rect 255635 297876 255636 297940
rect 255700 297876 255701 297940
rect 255635 297875 255701 297876
rect 256742 297805 256802 299782
rect 257064 299570 257124 300106
rect 257880 299570 257940 300106
rect 257064 299510 257170 299570
rect 257110 297941 257170 299510
rect 257846 299510 257940 299570
rect 258288 299570 258348 300106
rect 259104 299570 259164 300106
rect 259376 299570 259436 300106
rect 258288 299510 258458 299570
rect 259104 299510 259194 299570
rect 257846 298213 257906 299510
rect 257843 298212 257909 298213
rect 257843 298148 257844 298212
rect 257908 298148 257909 298212
rect 257843 298147 257909 298148
rect 257107 297940 257173 297941
rect 257107 297876 257108 297940
rect 257172 297876 257173 297940
rect 257107 297875 257173 297876
rect 256739 297804 256805 297805
rect 256739 297740 256740 297804
rect 256804 297740 256805 297804
rect 256739 297739 256805 297740
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 252000 254414 254898
rect 257514 295174 258134 298000
rect 258398 297805 258458 299510
rect 259134 297941 259194 299510
rect 259318 299510 259436 299570
rect 260600 299570 260660 300106
rect 260736 299570 260796 300106
rect 261416 299570 261476 300106
rect 261824 299570 261884 300106
rect 262912 299570 262972 300106
rect 263184 299570 263244 300106
rect 260600 299510 260666 299570
rect 260736 299510 260850 299570
rect 261416 299510 261586 299570
rect 261824 299510 261954 299570
rect 262912 299510 263058 299570
rect 259318 298077 259378 299510
rect 259315 298076 259381 298077
rect 259315 298012 259316 298076
rect 259380 298012 259381 298076
rect 259315 298011 259381 298012
rect 260606 297941 260666 299510
rect 260790 298077 260850 299510
rect 261526 298213 261586 299510
rect 261894 298213 261954 299510
rect 261523 298212 261589 298213
rect 261523 298148 261524 298212
rect 261588 298148 261589 298212
rect 261523 298147 261589 298148
rect 261891 298212 261957 298213
rect 261891 298148 261892 298212
rect 261956 298148 261957 298212
rect 261891 298147 261957 298148
rect 260787 298076 260853 298077
rect 260787 298012 260788 298076
rect 260852 298012 260853 298076
rect 260787 298011 260853 298012
rect 259131 297940 259197 297941
rect 259131 297876 259132 297940
rect 259196 297876 259197 297940
rect 259131 297875 259197 297876
rect 260603 297940 260669 297941
rect 260603 297876 260604 297940
rect 260668 297876 260669 297940
rect 260603 297875 260669 297876
rect 258395 297804 258461 297805
rect 258395 297740 258396 297804
rect 258460 297740 258461 297804
rect 258395 297739 258461 297740
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 252000 258134 258618
rect 261234 262894 261854 298000
rect 262998 297941 263058 299510
rect 263182 299510 263244 299570
rect 264000 299570 264060 300106
rect 264408 299570 264468 300106
rect 265224 299570 265284 300106
rect 264000 299510 264162 299570
rect 264408 299510 264530 299570
rect 263182 298077 263242 299510
rect 263179 298076 263245 298077
rect 263179 298012 263180 298076
rect 263244 298012 263245 298076
rect 263179 298011 263245 298012
rect 262995 297940 263061 297941
rect 262995 297876 262996 297940
rect 263060 297876 263061 297940
rect 262995 297875 263061 297876
rect 264102 296989 264162 299510
rect 264099 296988 264165 296989
rect 264099 296924 264100 296988
rect 264164 296924 264165 296988
rect 264099 296923 264165 296924
rect 264470 296853 264530 299510
rect 265206 299510 265284 299570
rect 265632 299570 265692 300106
rect 266584 299570 266644 300106
rect 266856 299570 266916 300106
rect 267672 299570 267732 300106
rect 265632 299510 265818 299570
rect 266584 299510 266738 299570
rect 266856 299510 266922 299570
rect 265206 298213 265266 299510
rect 265203 298212 265269 298213
rect 265203 298148 265204 298212
rect 265268 298148 265269 298212
rect 265203 298147 265269 298148
rect 264467 296852 264533 296853
rect 264467 296788 264468 296852
rect 264532 296788 264533 296852
rect 264467 296787 264533 296788
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 252000 261854 262338
rect 264954 266614 265574 298000
rect 265758 296853 265818 299510
rect 266678 296989 266738 299510
rect 266862 297125 266922 299510
rect 267598 299510 267732 299570
rect 267808 299570 267868 300106
rect 269304 299570 269364 300106
rect 267808 299510 268026 299570
rect 266859 297124 266925 297125
rect 266859 297060 266860 297124
rect 266924 297060 266925 297124
rect 266859 297059 266925 297060
rect 266675 296988 266741 296989
rect 266675 296924 266676 296988
rect 266740 296924 266741 296988
rect 266675 296923 266741 296924
rect 267598 296853 267658 299510
rect 267966 296853 268026 299510
rect 269254 299510 269364 299570
rect 270528 299570 270588 300106
rect 271888 299570 271948 300106
rect 270528 299510 270602 299570
rect 269254 296853 269314 299510
rect 270542 296853 270602 299510
rect 271830 299510 271948 299570
rect 273112 299570 273172 300106
rect 274336 299842 274396 300106
rect 274336 299782 274466 299842
rect 273112 299510 273178 299570
rect 271830 298213 271890 299510
rect 271827 298212 271893 298213
rect 271827 298148 271828 298212
rect 271892 298148 271893 298212
rect 271827 298147 271893 298148
rect 265755 296852 265821 296853
rect 265755 296788 265756 296852
rect 265820 296788 265821 296852
rect 265755 296787 265821 296788
rect 267595 296852 267661 296853
rect 267595 296788 267596 296852
rect 267660 296788 267661 296852
rect 267595 296787 267661 296788
rect 267963 296852 268029 296853
rect 267963 296788 267964 296852
rect 268028 296788 268029 296852
rect 267963 296787 268029 296788
rect 269251 296852 269317 296853
rect 269251 296788 269252 296852
rect 269316 296788 269317 296852
rect 269251 296787 269317 296788
rect 270539 296852 270605 296853
rect 270539 296788 270540 296852
rect 270604 296788 270605 296852
rect 270539 296787 270605 296788
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 252000 265574 266058
rect 271794 273454 272414 298000
rect 273118 296853 273178 299510
rect 274406 298077 274466 299782
rect 275560 299570 275620 300106
rect 275510 299510 275620 299570
rect 276784 299570 276844 300106
rect 276784 299510 276858 299570
rect 275510 298213 275570 299510
rect 275507 298212 275573 298213
rect 275507 298148 275508 298212
rect 275572 298148 275573 298212
rect 275507 298147 275573 298148
rect 276798 298077 276858 299510
rect 274403 298076 274469 298077
rect 274403 298012 274404 298076
rect 274468 298012 274469 298076
rect 274403 298011 274469 298012
rect 276795 298076 276861 298077
rect 276795 298012 276796 298076
rect 276860 298012 276861 298076
rect 276795 298011 276861 298012
rect 273115 296852 273181 296853
rect 273115 296788 273116 296852
rect 273180 296788 273181 296852
rect 273115 296787 273181 296788
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 252000 272414 272898
rect 275514 277174 276134 298000
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 252000 276134 276618
rect 279234 280894 279854 298000
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 252000 279854 280338
rect 282954 284614 283574 298000
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 252000 283574 284058
rect 289794 291454 290414 298000
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 252000 290414 254898
rect 293514 295174 294134 298000
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 252000 294134 258618
rect 297234 262894 297854 298000
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 252000 297854 262338
rect 300954 266614 301574 298000
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 252000 301574 266058
rect 307794 273454 308414 298000
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 252000 308414 272898
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 252000 312134 276618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 252000 315854 280338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 252000 319574 284058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 252000 326414 254898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 252000 330134 258618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 252000 333854 262338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 252000 337574 266058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 252000 344414 272898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 252000 348134 276618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 252000 351854 280338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 252000 355574 284058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 252000 362414 254898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 252000 366134 258618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 252000 369854 262338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 252000 373574 266058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 252000 380414 272898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 252000 384134 276618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 252000 387854 280338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 252000 391574 284058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 252000 398414 254898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 252000 402134 258618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408539 297532 408605 297533
rect 408539 297468 408540 297532
rect 408604 297468 408605 297532
rect 408539 297467 408605 297468
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 252000 405854 262338
rect 209568 237454 209888 237486
rect 209568 237218 209610 237454
rect 209846 237218 209888 237454
rect 209568 237134 209888 237218
rect 209568 236898 209610 237134
rect 209846 236898 209888 237134
rect 209568 236866 209888 236898
rect 240288 237454 240608 237486
rect 240288 237218 240330 237454
rect 240566 237218 240608 237454
rect 240288 237134 240608 237218
rect 240288 236898 240330 237134
rect 240566 236898 240608 237134
rect 240288 236866 240608 236898
rect 271008 237454 271328 237486
rect 271008 237218 271050 237454
rect 271286 237218 271328 237454
rect 271008 237134 271328 237218
rect 271008 236898 271050 237134
rect 271286 236898 271328 237134
rect 271008 236866 271328 236898
rect 301728 237454 302048 237486
rect 301728 237218 301770 237454
rect 302006 237218 302048 237454
rect 301728 237134 302048 237218
rect 301728 236898 301770 237134
rect 302006 236898 302048 237134
rect 301728 236866 302048 236898
rect 332448 237454 332768 237486
rect 332448 237218 332490 237454
rect 332726 237218 332768 237454
rect 332448 237134 332768 237218
rect 332448 236898 332490 237134
rect 332726 236898 332768 237134
rect 332448 236866 332768 236898
rect 363168 237454 363488 237486
rect 363168 237218 363210 237454
rect 363446 237218 363488 237454
rect 363168 237134 363488 237218
rect 363168 236898 363210 237134
rect 363446 236898 363488 237134
rect 363168 236866 363488 236898
rect 393888 237454 394208 237486
rect 393888 237218 393930 237454
rect 394166 237218 394208 237454
rect 393888 237134 394208 237218
rect 393888 236898 393930 237134
rect 394166 236898 394208 237134
rect 393888 236866 394208 236898
rect 408542 234290 408602 297467
rect 408723 297396 408789 297397
rect 408723 297332 408724 297396
rect 408788 297332 408789 297396
rect 408723 297331 408789 297332
rect 408726 238770 408786 297331
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 252000 409574 266058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 409275 251836 409341 251837
rect 409275 251772 409276 251836
rect 409340 251772 409341 251836
rect 409275 251771 409341 251772
rect 409278 248301 409338 251771
rect 409275 248300 409341 248301
rect 409275 248236 409276 248300
rect 409340 248236 409341 248300
rect 409275 248235 409341 248236
rect 408726 238710 409338 238770
rect 409278 237829 409338 238710
rect 409275 237828 409341 237829
rect 409275 237764 409276 237828
rect 409340 237764 409341 237828
rect 409275 237763 409341 237764
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 409275 234292 409341 234293
rect 409275 234290 409276 234292
rect 408542 234230 409276 234290
rect 409275 234228 409276 234230
rect 409340 234228 409341 234292
rect 409275 234227 409341 234228
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 194208 219454 194528 219486
rect 194208 219218 194250 219454
rect 194486 219218 194528 219454
rect 194208 219134 194528 219218
rect 194208 218898 194250 219134
rect 194486 218898 194528 219134
rect 194208 218866 194528 218898
rect 224928 219454 225248 219486
rect 224928 219218 224970 219454
rect 225206 219218 225248 219454
rect 224928 219134 225248 219218
rect 224928 218898 224970 219134
rect 225206 218898 225248 219134
rect 224928 218866 225248 218898
rect 255648 219454 255968 219486
rect 255648 219218 255690 219454
rect 255926 219218 255968 219454
rect 255648 219134 255968 219218
rect 255648 218898 255690 219134
rect 255926 218898 255968 219134
rect 255648 218866 255968 218898
rect 286368 219454 286688 219486
rect 286368 219218 286410 219454
rect 286646 219218 286688 219454
rect 286368 219134 286688 219218
rect 286368 218898 286410 219134
rect 286646 218898 286688 219134
rect 286368 218866 286688 218898
rect 317088 219454 317408 219486
rect 317088 219218 317130 219454
rect 317366 219218 317408 219454
rect 317088 219134 317408 219218
rect 317088 218898 317130 219134
rect 317366 218898 317408 219134
rect 317088 218866 317408 218898
rect 347808 219454 348128 219486
rect 347808 219218 347850 219454
rect 348086 219218 348128 219454
rect 347808 219134 348128 219218
rect 347808 218898 347850 219134
rect 348086 218898 348128 219134
rect 347808 218866 348128 218898
rect 378528 219454 378848 219486
rect 378528 219218 378570 219454
rect 378806 219218 378848 219454
rect 378528 219134 378848 219218
rect 378528 218898 378570 219134
rect 378806 218898 378848 219134
rect 378528 218866 378848 218898
rect 209568 201454 209888 201486
rect 209568 201218 209610 201454
rect 209846 201218 209888 201454
rect 209568 201134 209888 201218
rect 209568 200898 209610 201134
rect 209846 200898 209888 201134
rect 209568 200866 209888 200898
rect 240288 201454 240608 201486
rect 240288 201218 240330 201454
rect 240566 201218 240608 201454
rect 240288 201134 240608 201218
rect 240288 200898 240330 201134
rect 240566 200898 240608 201134
rect 240288 200866 240608 200898
rect 271008 201454 271328 201486
rect 271008 201218 271050 201454
rect 271286 201218 271328 201454
rect 271008 201134 271328 201218
rect 271008 200898 271050 201134
rect 271286 200898 271328 201134
rect 271008 200866 271328 200898
rect 301728 201454 302048 201486
rect 301728 201218 301770 201454
rect 302006 201218 302048 201454
rect 301728 201134 302048 201218
rect 301728 200898 301770 201134
rect 302006 200898 302048 201134
rect 301728 200866 302048 200898
rect 332448 201454 332768 201486
rect 332448 201218 332490 201454
rect 332726 201218 332768 201454
rect 332448 201134 332768 201218
rect 332448 200898 332490 201134
rect 332726 200898 332768 201134
rect 332448 200866 332768 200898
rect 363168 201454 363488 201486
rect 363168 201218 363210 201454
rect 363446 201218 363488 201454
rect 363168 201134 363488 201218
rect 363168 200898 363210 201134
rect 363446 200898 363488 201134
rect 363168 200866 363488 200898
rect 393888 201454 394208 201486
rect 393888 201218 393930 201454
rect 394166 201218 394208 201454
rect 393888 201134 394208 201218
rect 393888 200898 393930 201134
rect 394166 200898 394208 201134
rect 393888 200866 394208 200898
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 194208 183454 194528 183486
rect 194208 183218 194250 183454
rect 194486 183218 194528 183454
rect 194208 183134 194528 183218
rect 194208 182898 194250 183134
rect 194486 182898 194528 183134
rect 194208 182866 194528 182898
rect 224928 183454 225248 183486
rect 224928 183218 224970 183454
rect 225206 183218 225248 183454
rect 224928 183134 225248 183218
rect 224928 182898 224970 183134
rect 225206 182898 225248 183134
rect 224928 182866 225248 182898
rect 255648 183454 255968 183486
rect 255648 183218 255690 183454
rect 255926 183218 255968 183454
rect 255648 183134 255968 183218
rect 255648 182898 255690 183134
rect 255926 182898 255968 183134
rect 255648 182866 255968 182898
rect 286368 183454 286688 183486
rect 286368 183218 286410 183454
rect 286646 183218 286688 183454
rect 286368 183134 286688 183218
rect 286368 182898 286410 183134
rect 286646 182898 286688 183134
rect 286368 182866 286688 182898
rect 317088 183454 317408 183486
rect 317088 183218 317130 183454
rect 317366 183218 317408 183454
rect 317088 183134 317408 183218
rect 317088 182898 317130 183134
rect 317366 182898 317408 183134
rect 317088 182866 317408 182898
rect 347808 183454 348128 183486
rect 347808 183218 347850 183454
rect 348086 183218 348128 183454
rect 347808 183134 348128 183218
rect 347808 182898 347850 183134
rect 348086 182898 348128 183134
rect 347808 182866 348128 182898
rect 378528 183454 378848 183486
rect 378528 183218 378570 183454
rect 378806 183218 378848 183454
rect 378528 183134 378848 183218
rect 378528 182898 378570 183134
rect 378806 182898 378848 183134
rect 378528 182866 378848 182898
rect 209568 165454 209888 165486
rect 209568 165218 209610 165454
rect 209846 165218 209888 165454
rect 209568 165134 209888 165218
rect 209568 164898 209610 165134
rect 209846 164898 209888 165134
rect 209568 164866 209888 164898
rect 240288 165454 240608 165486
rect 240288 165218 240330 165454
rect 240566 165218 240608 165454
rect 240288 165134 240608 165218
rect 240288 164898 240330 165134
rect 240566 164898 240608 165134
rect 240288 164866 240608 164898
rect 271008 165454 271328 165486
rect 271008 165218 271050 165454
rect 271286 165218 271328 165454
rect 271008 165134 271328 165218
rect 271008 164898 271050 165134
rect 271286 164898 271328 165134
rect 271008 164866 271328 164898
rect 301728 165454 302048 165486
rect 301728 165218 301770 165454
rect 302006 165218 302048 165454
rect 301728 165134 302048 165218
rect 301728 164898 301770 165134
rect 302006 164898 302048 165134
rect 301728 164866 302048 164898
rect 332448 165454 332768 165486
rect 332448 165218 332490 165454
rect 332726 165218 332768 165454
rect 332448 165134 332768 165218
rect 332448 164898 332490 165134
rect 332726 164898 332768 165134
rect 332448 164866 332768 164898
rect 363168 165454 363488 165486
rect 363168 165218 363210 165454
rect 363446 165218 363488 165454
rect 363168 165134 363488 165218
rect 363168 164898 363210 165134
rect 363446 164898 363488 165134
rect 363168 164866 363488 164898
rect 393888 165454 394208 165486
rect 393888 165218 393930 165454
rect 394166 165218 394208 165454
rect 393888 165134 394208 165218
rect 393888 164898 393930 165134
rect 394166 164898 394208 165134
rect 393888 164866 394208 164898
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 194208 147454 194528 147486
rect 194208 147218 194250 147454
rect 194486 147218 194528 147454
rect 194208 147134 194528 147218
rect 194208 146898 194250 147134
rect 194486 146898 194528 147134
rect 194208 146866 194528 146898
rect 224928 147454 225248 147486
rect 224928 147218 224970 147454
rect 225206 147218 225248 147454
rect 224928 147134 225248 147218
rect 224928 146898 224970 147134
rect 225206 146898 225248 147134
rect 224928 146866 225248 146898
rect 255648 147454 255968 147486
rect 255648 147218 255690 147454
rect 255926 147218 255968 147454
rect 255648 147134 255968 147218
rect 255648 146898 255690 147134
rect 255926 146898 255968 147134
rect 255648 146866 255968 146898
rect 286368 147454 286688 147486
rect 286368 147218 286410 147454
rect 286646 147218 286688 147454
rect 286368 147134 286688 147218
rect 286368 146898 286410 147134
rect 286646 146898 286688 147134
rect 286368 146866 286688 146898
rect 317088 147454 317408 147486
rect 317088 147218 317130 147454
rect 317366 147218 317408 147454
rect 317088 147134 317408 147218
rect 317088 146898 317130 147134
rect 317366 146898 317408 147134
rect 317088 146866 317408 146898
rect 347808 147454 348128 147486
rect 347808 147218 347850 147454
rect 348086 147218 348128 147454
rect 347808 147134 348128 147218
rect 347808 146898 347850 147134
rect 348086 146898 348128 147134
rect 347808 146866 348128 146898
rect 378528 147454 378848 147486
rect 378528 147218 378570 147454
rect 378806 147218 378848 147454
rect 378528 147134 378848 147218
rect 378528 146898 378570 147134
rect 378806 146898 378848 147134
rect 378528 146866 378848 146898
rect 209568 129454 209888 129486
rect 209568 129218 209610 129454
rect 209846 129218 209888 129454
rect 209568 129134 209888 129218
rect 209568 128898 209610 129134
rect 209846 128898 209888 129134
rect 209568 128866 209888 128898
rect 240288 129454 240608 129486
rect 240288 129218 240330 129454
rect 240566 129218 240608 129454
rect 240288 129134 240608 129218
rect 240288 128898 240330 129134
rect 240566 128898 240608 129134
rect 240288 128866 240608 128898
rect 271008 129454 271328 129486
rect 271008 129218 271050 129454
rect 271286 129218 271328 129454
rect 271008 129134 271328 129218
rect 271008 128898 271050 129134
rect 271286 128898 271328 129134
rect 271008 128866 271328 128898
rect 301728 129454 302048 129486
rect 301728 129218 301770 129454
rect 302006 129218 302048 129454
rect 301728 129134 302048 129218
rect 301728 128898 301770 129134
rect 302006 128898 302048 129134
rect 301728 128866 302048 128898
rect 332448 129454 332768 129486
rect 332448 129218 332490 129454
rect 332726 129218 332768 129454
rect 332448 129134 332768 129218
rect 332448 128898 332490 129134
rect 332726 128898 332768 129134
rect 332448 128866 332768 128898
rect 363168 129454 363488 129486
rect 363168 129218 363210 129454
rect 363446 129218 363488 129454
rect 363168 129134 363488 129218
rect 363168 128898 363210 129134
rect 363446 128898 363488 129134
rect 363168 128866 363488 128898
rect 393888 129454 394208 129486
rect 393888 129218 393930 129454
rect 394166 129218 394208 129454
rect 393888 129134 394208 129218
rect 393888 128898 393930 129134
rect 394166 128898 394208 129134
rect 393888 128866 394208 128898
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 194208 111454 194528 111486
rect 194208 111218 194250 111454
rect 194486 111218 194528 111454
rect 194208 111134 194528 111218
rect 194208 110898 194250 111134
rect 194486 110898 194528 111134
rect 194208 110866 194528 110898
rect 224928 111454 225248 111486
rect 224928 111218 224970 111454
rect 225206 111218 225248 111454
rect 224928 111134 225248 111218
rect 224928 110898 224970 111134
rect 225206 110898 225248 111134
rect 224928 110866 225248 110898
rect 255648 111454 255968 111486
rect 255648 111218 255690 111454
rect 255926 111218 255968 111454
rect 255648 111134 255968 111218
rect 255648 110898 255690 111134
rect 255926 110898 255968 111134
rect 255648 110866 255968 110898
rect 286368 111454 286688 111486
rect 286368 111218 286410 111454
rect 286646 111218 286688 111454
rect 286368 111134 286688 111218
rect 286368 110898 286410 111134
rect 286646 110898 286688 111134
rect 286368 110866 286688 110898
rect 317088 111454 317408 111486
rect 317088 111218 317130 111454
rect 317366 111218 317408 111454
rect 317088 111134 317408 111218
rect 317088 110898 317130 111134
rect 317366 110898 317408 111134
rect 317088 110866 317408 110898
rect 347808 111454 348128 111486
rect 347808 111218 347850 111454
rect 348086 111218 348128 111454
rect 347808 111134 348128 111218
rect 347808 110898 347850 111134
rect 348086 110898 348128 111134
rect 347808 110866 348128 110898
rect 378528 111454 378848 111486
rect 378528 111218 378570 111454
rect 378806 111218 378848 111454
rect 378528 111134 378848 111218
rect 378528 110898 378570 111134
rect 378806 110898 378848 111134
rect 378528 110866 378848 110898
rect 209568 93454 209888 93486
rect 209568 93218 209610 93454
rect 209846 93218 209888 93454
rect 209568 93134 209888 93218
rect 209568 92898 209610 93134
rect 209846 92898 209888 93134
rect 209568 92866 209888 92898
rect 240288 93454 240608 93486
rect 240288 93218 240330 93454
rect 240566 93218 240608 93454
rect 240288 93134 240608 93218
rect 240288 92898 240330 93134
rect 240566 92898 240608 93134
rect 240288 92866 240608 92898
rect 271008 93454 271328 93486
rect 271008 93218 271050 93454
rect 271286 93218 271328 93454
rect 271008 93134 271328 93218
rect 271008 92898 271050 93134
rect 271286 92898 271328 93134
rect 271008 92866 271328 92898
rect 301728 93454 302048 93486
rect 301728 93218 301770 93454
rect 302006 93218 302048 93454
rect 301728 93134 302048 93218
rect 301728 92898 301770 93134
rect 302006 92898 302048 93134
rect 301728 92866 302048 92898
rect 332448 93454 332768 93486
rect 332448 93218 332490 93454
rect 332726 93218 332768 93454
rect 332448 93134 332768 93218
rect 332448 92898 332490 93134
rect 332726 92898 332768 93134
rect 332448 92866 332768 92898
rect 363168 93454 363488 93486
rect 363168 93218 363210 93454
rect 363446 93218 363488 93454
rect 363168 93134 363488 93218
rect 363168 92898 363210 93134
rect 363446 92898 363488 93134
rect 363168 92866 363488 92898
rect 393888 93454 394208 93486
rect 393888 93218 393930 93454
rect 394166 93218 394208 93454
rect 393888 93134 394208 93218
rect 393888 92898 393930 93134
rect 394166 92898 394208 93134
rect 393888 92866 394208 92898
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 194208 75454 194528 75486
rect 194208 75218 194250 75454
rect 194486 75218 194528 75454
rect 194208 75134 194528 75218
rect 194208 74898 194250 75134
rect 194486 74898 194528 75134
rect 194208 74866 194528 74898
rect 224928 75454 225248 75486
rect 224928 75218 224970 75454
rect 225206 75218 225248 75454
rect 224928 75134 225248 75218
rect 224928 74898 224970 75134
rect 225206 74898 225248 75134
rect 224928 74866 225248 74898
rect 255648 75454 255968 75486
rect 255648 75218 255690 75454
rect 255926 75218 255968 75454
rect 255648 75134 255968 75218
rect 255648 74898 255690 75134
rect 255926 74898 255968 75134
rect 255648 74866 255968 74898
rect 286368 75454 286688 75486
rect 286368 75218 286410 75454
rect 286646 75218 286688 75454
rect 286368 75134 286688 75218
rect 286368 74898 286410 75134
rect 286646 74898 286688 75134
rect 286368 74866 286688 74898
rect 317088 75454 317408 75486
rect 317088 75218 317130 75454
rect 317366 75218 317408 75454
rect 317088 75134 317408 75218
rect 317088 74898 317130 75134
rect 317366 74898 317408 75134
rect 317088 74866 317408 74898
rect 347808 75454 348128 75486
rect 347808 75218 347850 75454
rect 348086 75218 348128 75454
rect 347808 75134 348128 75218
rect 347808 74898 347850 75134
rect 348086 74898 348128 75134
rect 347808 74866 348128 74898
rect 378528 75454 378848 75486
rect 378528 75218 378570 75454
rect 378806 75218 378848 75454
rect 378528 75134 378848 75218
rect 378528 74898 378570 75134
rect 378806 74898 378848 75134
rect 378528 74866 378848 74898
rect 209568 57454 209888 57486
rect 209568 57218 209610 57454
rect 209846 57218 209888 57454
rect 209568 57134 209888 57218
rect 209568 56898 209610 57134
rect 209846 56898 209888 57134
rect 209568 56866 209888 56898
rect 240288 57454 240608 57486
rect 240288 57218 240330 57454
rect 240566 57218 240608 57454
rect 240288 57134 240608 57218
rect 240288 56898 240330 57134
rect 240566 56898 240608 57134
rect 240288 56866 240608 56898
rect 271008 57454 271328 57486
rect 271008 57218 271050 57454
rect 271286 57218 271328 57454
rect 271008 57134 271328 57218
rect 271008 56898 271050 57134
rect 271286 56898 271328 57134
rect 271008 56866 271328 56898
rect 301728 57454 302048 57486
rect 301728 57218 301770 57454
rect 302006 57218 302048 57454
rect 301728 57134 302048 57218
rect 301728 56898 301770 57134
rect 302006 56898 302048 57134
rect 301728 56866 302048 56898
rect 332448 57454 332768 57486
rect 332448 57218 332490 57454
rect 332726 57218 332768 57454
rect 332448 57134 332768 57218
rect 332448 56898 332490 57134
rect 332726 56898 332768 57134
rect 332448 56866 332768 56898
rect 363168 57454 363488 57486
rect 363168 57218 363210 57454
rect 363446 57218 363488 57454
rect 363168 57134 363488 57218
rect 363168 56898 363210 57134
rect 363446 56898 363488 57134
rect 363168 56866 363488 56898
rect 393888 57454 394208 57486
rect 393888 57218 393930 57454
rect 394166 57218 394208 57454
rect 393888 57134 394208 57218
rect 393888 56898 393930 57134
rect 394166 56898 394208 57134
rect 393888 56866 394208 56898
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 194208 39454 194528 39486
rect 194208 39218 194250 39454
rect 194486 39218 194528 39454
rect 194208 39134 194528 39218
rect 194208 38898 194250 39134
rect 194486 38898 194528 39134
rect 194208 38866 194528 38898
rect 224928 39454 225248 39486
rect 224928 39218 224970 39454
rect 225206 39218 225248 39454
rect 224928 39134 225248 39218
rect 224928 38898 224970 39134
rect 225206 38898 225248 39134
rect 224928 38866 225248 38898
rect 255648 39454 255968 39486
rect 255648 39218 255690 39454
rect 255926 39218 255968 39454
rect 255648 39134 255968 39218
rect 255648 38898 255690 39134
rect 255926 38898 255968 39134
rect 255648 38866 255968 38898
rect 286368 39454 286688 39486
rect 286368 39218 286410 39454
rect 286646 39218 286688 39454
rect 286368 39134 286688 39218
rect 286368 38898 286410 39134
rect 286646 38898 286688 39134
rect 286368 38866 286688 38898
rect 317088 39454 317408 39486
rect 317088 39218 317130 39454
rect 317366 39218 317408 39454
rect 317088 39134 317408 39218
rect 317088 38898 317130 39134
rect 317366 38898 317408 39134
rect 317088 38866 317408 38898
rect 347808 39454 348128 39486
rect 347808 39218 347850 39454
rect 348086 39218 348128 39454
rect 347808 39134 348128 39218
rect 347808 38898 347850 39134
rect 348086 38898 348128 39134
rect 347808 38866 348128 38898
rect 378528 39454 378848 39486
rect 378528 39218 378570 39454
rect 378806 39218 378848 39454
rect 378528 39134 378848 39218
rect 378528 38898 378570 39134
rect 378806 38898 378848 39134
rect 378528 38866 378848 38898
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 28000
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 28000
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 28000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 28000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 28000
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 28000
rect 217794 3454 218414 28000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 7174 222134 28000
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 10894 225854 28000
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 28000
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 28000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 28000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 28000
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 28000
rect 253794 3454 254414 28000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 28000
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 28000
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 28000
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 28000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 28000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 28000
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 28000
rect 289794 3454 290414 28000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 7174 294134 28000
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 10894 297854 28000
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 28000
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 21454 308414 28000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 28000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 -5146 315854 28000
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 28000
rect 325794 3454 326414 28000
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 7174 330134 28000
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 10894 333854 28000
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 14614 337574 28000
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 21454 344414 28000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 28000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 -5146 351854 28000
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 28000
rect 361794 3454 362414 28000
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 7174 366134 28000
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 10894 369854 28000
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 14614 373574 28000
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 28000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 28000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 -5146 387854 28000
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 28000
rect 397794 3454 398414 28000
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 7174 402134 28000
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 10894 405854 28000
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 14614 409574 28000
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 132000 438134 150618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 132000 441854 154338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 132000 445574 158058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 132000 452414 164898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 132000 456134 132618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 132000 459854 136338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 132000 463574 140058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 132000 470414 146898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 132000 474134 150618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 132000 477854 154338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 132000 481574 158058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 132000 488414 164898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 132000 492134 132618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 132000 495854 136338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 132000 499574 140058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 132000 506414 146898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 132000 510134 150618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 132000 513854 154338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 132000 517574 158058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 132000 524414 164898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 132000 528134 132618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 132000 531854 136338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 132000 535574 140058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 132000 542414 146898
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 444208 111454 444528 111486
rect 444208 111218 444250 111454
rect 444486 111218 444528 111454
rect 444208 111134 444528 111218
rect 444208 110898 444250 111134
rect 444486 110898 444528 111134
rect 444208 110866 444528 110898
rect 474928 111454 475248 111486
rect 474928 111218 474970 111454
rect 475206 111218 475248 111454
rect 474928 111134 475248 111218
rect 474928 110898 474970 111134
rect 475206 110898 475248 111134
rect 474928 110866 475248 110898
rect 505648 111454 505968 111486
rect 505648 111218 505690 111454
rect 505926 111218 505968 111454
rect 505648 111134 505968 111218
rect 505648 110898 505690 111134
rect 505926 110898 505968 111134
rect 505648 110866 505968 110898
rect 536368 111454 536688 111486
rect 536368 111218 536410 111454
rect 536646 111218 536688 111454
rect 536368 111134 536688 111218
rect 536368 110898 536410 111134
rect 536646 110898 536688 111134
rect 536368 110866 536688 110898
rect 459568 93454 459888 93486
rect 459568 93218 459610 93454
rect 459846 93218 459888 93454
rect 459568 93134 459888 93218
rect 459568 92898 459610 93134
rect 459846 92898 459888 93134
rect 459568 92866 459888 92898
rect 490288 93454 490608 93486
rect 490288 93218 490330 93454
rect 490566 93218 490608 93454
rect 490288 93134 490608 93218
rect 490288 92898 490330 93134
rect 490566 92898 490608 93134
rect 490288 92866 490608 92898
rect 521008 93454 521328 93486
rect 521008 93218 521050 93454
rect 521286 93218 521328 93454
rect 521008 93134 521328 93218
rect 521008 92898 521050 93134
rect 521286 92898 521328 93134
rect 521008 92866 521328 92898
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 444208 75454 444528 75486
rect 444208 75218 444250 75454
rect 444486 75218 444528 75454
rect 444208 75134 444528 75218
rect 444208 74898 444250 75134
rect 444486 74898 444528 75134
rect 444208 74866 444528 74898
rect 474928 75454 475248 75486
rect 474928 75218 474970 75454
rect 475206 75218 475248 75454
rect 474928 75134 475248 75218
rect 474928 74898 474970 75134
rect 475206 74898 475248 75134
rect 474928 74866 475248 74898
rect 505648 75454 505968 75486
rect 505648 75218 505690 75454
rect 505926 75218 505968 75454
rect 505648 75134 505968 75218
rect 505648 74898 505690 75134
rect 505926 74898 505968 75134
rect 505648 74866 505968 74898
rect 536368 75454 536688 75486
rect 536368 75218 536410 75454
rect 536646 75218 536688 75454
rect 536368 75134 536688 75218
rect 536368 74898 536410 75134
rect 536646 74898 536688 75134
rect 536368 74866 536688 74898
rect 459568 57454 459888 57486
rect 459568 57218 459610 57454
rect 459846 57218 459888 57454
rect 459568 57134 459888 57218
rect 459568 56898 459610 57134
rect 459846 56898 459888 57134
rect 459568 56866 459888 56898
rect 490288 57454 490608 57486
rect 490288 57218 490330 57454
rect 490566 57218 490608 57454
rect 490288 57134 490608 57218
rect 490288 56898 490330 57134
rect 490566 56898 490608 57134
rect 490288 56866 490608 56898
rect 521008 57454 521328 57486
rect 521008 57218 521050 57454
rect 521286 57218 521328 57454
rect 521008 57134 521328 57218
rect 521008 56898 521050 57134
rect 521286 56898 521328 57134
rect 521008 56866 521328 56898
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 444208 39454 444528 39486
rect 444208 39218 444250 39454
rect 444486 39218 444528 39454
rect 444208 39134 444528 39218
rect 444208 38898 444250 39134
rect 444486 38898 444528 39134
rect 444208 38866 444528 38898
rect 474928 39454 475248 39486
rect 474928 39218 474970 39454
rect 475206 39218 475248 39454
rect 474928 39134 475248 39218
rect 474928 38898 474970 39134
rect 475206 38898 475248 39134
rect 474928 38866 475248 38898
rect 505648 39454 505968 39486
rect 505648 39218 505690 39454
rect 505926 39218 505968 39454
rect 505648 39134 505968 39218
rect 505648 38898 505690 39134
rect 505926 38898 505968 39134
rect 505648 38866 505968 38898
rect 536368 39454 536688 39486
rect 536368 39218 536410 39454
rect 536646 39218 536688 39454
rect 536368 39134 536688 39218
rect 536368 38898 536410 39134
rect 536646 38898 536688 39134
rect 536368 38866 536688 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 7174 438134 28000
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 10894 441854 28000
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 14614 445574 28000
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 21454 452414 28000
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 28000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 -5146 459854 28000
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 28000
rect 469794 3454 470414 28000
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 7174 474134 28000
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 10894 477854 28000
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 14614 481574 28000
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 21454 488414 28000
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 28000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 -5146 495854 28000
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 28000
rect 505794 3454 506414 28000
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 7174 510134 28000
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 10894 513854 28000
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 14614 517574 28000
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 21454 524414 28000
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 25174 528134 28000
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 -5146 531854 28000
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 28000
rect 541794 3454 542414 28000
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 51008 363218 51244 363454
rect 51008 362898 51244 363134
rect 144712 363218 144948 363454
rect 144712 362898 144948 363134
rect 50328 345218 50564 345454
rect 50328 344898 50564 345134
rect 145392 345218 145628 345454
rect 145392 344898 145628 345134
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 51008 327218 51244 327454
rect 51008 326898 51244 327134
rect 144712 327218 144948 327454
rect 144712 326898 144948 327134
rect 50328 309218 50564 309454
rect 50328 308898 50564 309134
rect 145392 309218 145628 309454
rect 145392 308898 145628 309134
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 34250 111218 34486 111454
rect 34250 110898 34486 111134
rect 64970 111218 65206 111454
rect 64970 110898 65206 111134
rect 95690 111218 95926 111454
rect 95690 110898 95926 111134
rect 126410 111218 126646 111454
rect 126410 110898 126646 111134
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 49610 93218 49846 93454
rect 49610 92898 49846 93134
rect 80330 93218 80566 93454
rect 80330 92898 80566 93134
rect 111050 93218 111286 93454
rect 111050 92898 111286 93134
rect 34250 75218 34486 75454
rect 34250 74898 34486 75134
rect 64970 75218 65206 75454
rect 64970 74898 65206 75134
rect 95690 75218 95926 75454
rect 95690 74898 95926 75134
rect 126410 75218 126646 75454
rect 126410 74898 126646 75134
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 49610 57218 49846 57454
rect 49610 56898 49846 57134
rect 80330 57218 80566 57454
rect 80330 56898 80566 57134
rect 111050 57218 111286 57454
rect 111050 56898 111286 57134
rect 34250 39218 34486 39454
rect 34250 38898 34486 39134
rect 64970 39218 65206 39454
rect 64970 38898 65206 39134
rect 95690 39218 95926 39454
rect 95690 38898 95926 39134
rect 126410 39218 126646 39454
rect 126410 38898 126646 39134
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 211008 363218 211244 363454
rect 211008 362898 211244 363134
rect 304712 363218 304948 363454
rect 304712 362898 304948 363134
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 210328 345218 210564 345454
rect 210328 344898 210564 345134
rect 305392 345218 305628 345454
rect 305392 344898 305628 345134
rect 211008 327218 211244 327454
rect 211008 326898 211244 327134
rect 304712 327218 304948 327454
rect 304712 326898 304948 327134
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 210328 309218 210564 309454
rect 210328 308898 210564 309134
rect 305392 309218 305628 309454
rect 305392 308898 305628 309134
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 209610 237218 209846 237454
rect 209610 236898 209846 237134
rect 240330 237218 240566 237454
rect 240330 236898 240566 237134
rect 271050 237218 271286 237454
rect 271050 236898 271286 237134
rect 301770 237218 302006 237454
rect 301770 236898 302006 237134
rect 332490 237218 332726 237454
rect 332490 236898 332726 237134
rect 363210 237218 363446 237454
rect 363210 236898 363446 237134
rect 393930 237218 394166 237454
rect 393930 236898 394166 237134
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 194250 219218 194486 219454
rect 194250 218898 194486 219134
rect 224970 219218 225206 219454
rect 224970 218898 225206 219134
rect 255690 219218 255926 219454
rect 255690 218898 255926 219134
rect 286410 219218 286646 219454
rect 286410 218898 286646 219134
rect 317130 219218 317366 219454
rect 317130 218898 317366 219134
rect 347850 219218 348086 219454
rect 347850 218898 348086 219134
rect 378570 219218 378806 219454
rect 378570 218898 378806 219134
rect 209610 201218 209846 201454
rect 209610 200898 209846 201134
rect 240330 201218 240566 201454
rect 240330 200898 240566 201134
rect 271050 201218 271286 201454
rect 271050 200898 271286 201134
rect 301770 201218 302006 201454
rect 301770 200898 302006 201134
rect 332490 201218 332726 201454
rect 332490 200898 332726 201134
rect 363210 201218 363446 201454
rect 363210 200898 363446 201134
rect 393930 201218 394166 201454
rect 393930 200898 394166 201134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 194250 183218 194486 183454
rect 194250 182898 194486 183134
rect 224970 183218 225206 183454
rect 224970 182898 225206 183134
rect 255690 183218 255926 183454
rect 255690 182898 255926 183134
rect 286410 183218 286646 183454
rect 286410 182898 286646 183134
rect 317130 183218 317366 183454
rect 317130 182898 317366 183134
rect 347850 183218 348086 183454
rect 347850 182898 348086 183134
rect 378570 183218 378806 183454
rect 378570 182898 378806 183134
rect 209610 165218 209846 165454
rect 209610 164898 209846 165134
rect 240330 165218 240566 165454
rect 240330 164898 240566 165134
rect 271050 165218 271286 165454
rect 271050 164898 271286 165134
rect 301770 165218 302006 165454
rect 301770 164898 302006 165134
rect 332490 165218 332726 165454
rect 332490 164898 332726 165134
rect 363210 165218 363446 165454
rect 363210 164898 363446 165134
rect 393930 165218 394166 165454
rect 393930 164898 394166 165134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 194250 147218 194486 147454
rect 194250 146898 194486 147134
rect 224970 147218 225206 147454
rect 224970 146898 225206 147134
rect 255690 147218 255926 147454
rect 255690 146898 255926 147134
rect 286410 147218 286646 147454
rect 286410 146898 286646 147134
rect 317130 147218 317366 147454
rect 317130 146898 317366 147134
rect 347850 147218 348086 147454
rect 347850 146898 348086 147134
rect 378570 147218 378806 147454
rect 378570 146898 378806 147134
rect 209610 129218 209846 129454
rect 209610 128898 209846 129134
rect 240330 129218 240566 129454
rect 240330 128898 240566 129134
rect 271050 129218 271286 129454
rect 271050 128898 271286 129134
rect 301770 129218 302006 129454
rect 301770 128898 302006 129134
rect 332490 129218 332726 129454
rect 332490 128898 332726 129134
rect 363210 129218 363446 129454
rect 363210 128898 363446 129134
rect 393930 129218 394166 129454
rect 393930 128898 394166 129134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 194250 111218 194486 111454
rect 194250 110898 194486 111134
rect 224970 111218 225206 111454
rect 224970 110898 225206 111134
rect 255690 111218 255926 111454
rect 255690 110898 255926 111134
rect 286410 111218 286646 111454
rect 286410 110898 286646 111134
rect 317130 111218 317366 111454
rect 317130 110898 317366 111134
rect 347850 111218 348086 111454
rect 347850 110898 348086 111134
rect 378570 111218 378806 111454
rect 378570 110898 378806 111134
rect 209610 93218 209846 93454
rect 209610 92898 209846 93134
rect 240330 93218 240566 93454
rect 240330 92898 240566 93134
rect 271050 93218 271286 93454
rect 271050 92898 271286 93134
rect 301770 93218 302006 93454
rect 301770 92898 302006 93134
rect 332490 93218 332726 93454
rect 332490 92898 332726 93134
rect 363210 93218 363446 93454
rect 363210 92898 363446 93134
rect 393930 93218 394166 93454
rect 393930 92898 394166 93134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 194250 75218 194486 75454
rect 194250 74898 194486 75134
rect 224970 75218 225206 75454
rect 224970 74898 225206 75134
rect 255690 75218 255926 75454
rect 255690 74898 255926 75134
rect 286410 75218 286646 75454
rect 286410 74898 286646 75134
rect 317130 75218 317366 75454
rect 317130 74898 317366 75134
rect 347850 75218 348086 75454
rect 347850 74898 348086 75134
rect 378570 75218 378806 75454
rect 378570 74898 378806 75134
rect 209610 57218 209846 57454
rect 209610 56898 209846 57134
rect 240330 57218 240566 57454
rect 240330 56898 240566 57134
rect 271050 57218 271286 57454
rect 271050 56898 271286 57134
rect 301770 57218 302006 57454
rect 301770 56898 302006 57134
rect 332490 57218 332726 57454
rect 332490 56898 332726 57134
rect 363210 57218 363446 57454
rect 363210 56898 363446 57134
rect 393930 57218 394166 57454
rect 393930 56898 394166 57134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 194250 39218 194486 39454
rect 194250 38898 194486 39134
rect 224970 39218 225206 39454
rect 224970 38898 225206 39134
rect 255690 39218 255926 39454
rect 255690 38898 255926 39134
rect 286410 39218 286646 39454
rect 286410 38898 286646 39134
rect 317130 39218 317366 39454
rect 317130 38898 317366 39134
rect 347850 39218 348086 39454
rect 347850 38898 348086 39134
rect 378570 39218 378806 39454
rect 378570 38898 378806 39134
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 444250 111218 444486 111454
rect 444250 110898 444486 111134
rect 474970 111218 475206 111454
rect 474970 110898 475206 111134
rect 505690 111218 505926 111454
rect 505690 110898 505926 111134
rect 536410 111218 536646 111454
rect 536410 110898 536646 111134
rect 459610 93218 459846 93454
rect 459610 92898 459846 93134
rect 490330 93218 490566 93454
rect 490330 92898 490566 93134
rect 521050 93218 521286 93454
rect 521050 92898 521286 93134
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 444250 75218 444486 75454
rect 444250 74898 444486 75134
rect 474970 75218 475206 75454
rect 474970 74898 475206 75134
rect 505690 75218 505926 75454
rect 505690 74898 505926 75134
rect 536410 75218 536646 75454
rect 536410 74898 536646 75134
rect 459610 57218 459846 57454
rect 459610 56898 459846 57134
rect 490330 57218 490566 57454
rect 490330 56898 490566 57134
rect 521050 57218 521286 57454
rect 521050 56898 521286 57134
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 444250 39218 444486 39454
rect 444250 38898 444486 39134
rect 474970 39218 475206 39454
rect 474970 38898 475206 39134
rect 505690 39218 505926 39454
rect 505690 38898 505926 39134
rect 536410 39218 536646 39454
rect 536410 38898 536646 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 51008 363454
rect 51244 363218 144712 363454
rect 144948 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 211008 363454
rect 211244 363218 304712 363454
rect 304948 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 51008 363134
rect 51244 362898 144712 363134
rect 144948 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 211008 363134
rect 211244 362898 304712 363134
rect 304948 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 50328 345454
rect 50564 345218 145392 345454
rect 145628 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 210328 345454
rect 210564 345218 305392 345454
rect 305628 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 50328 345134
rect 50564 344898 145392 345134
rect 145628 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 210328 345134
rect 210564 344898 305392 345134
rect 305628 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 51008 327454
rect 51244 327218 144712 327454
rect 144948 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 211008 327454
rect 211244 327218 304712 327454
rect 304948 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 51008 327134
rect 51244 326898 144712 327134
rect 144948 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 211008 327134
rect 211244 326898 304712 327134
rect 304948 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 50328 309454
rect 50564 309218 145392 309454
rect 145628 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 210328 309454
rect 210564 309218 305392 309454
rect 305628 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 50328 309134
rect 50564 308898 145392 309134
rect 145628 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 210328 309134
rect 210564 308898 305392 309134
rect 305628 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 209610 237454
rect 209846 237218 240330 237454
rect 240566 237218 271050 237454
rect 271286 237218 301770 237454
rect 302006 237218 332490 237454
rect 332726 237218 363210 237454
rect 363446 237218 393930 237454
rect 394166 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 209610 237134
rect 209846 236898 240330 237134
rect 240566 236898 271050 237134
rect 271286 236898 301770 237134
rect 302006 236898 332490 237134
rect 332726 236898 363210 237134
rect 363446 236898 393930 237134
rect 394166 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 194250 219454
rect 194486 219218 224970 219454
rect 225206 219218 255690 219454
rect 255926 219218 286410 219454
rect 286646 219218 317130 219454
rect 317366 219218 347850 219454
rect 348086 219218 378570 219454
rect 378806 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 194250 219134
rect 194486 218898 224970 219134
rect 225206 218898 255690 219134
rect 255926 218898 286410 219134
rect 286646 218898 317130 219134
rect 317366 218898 347850 219134
rect 348086 218898 378570 219134
rect 378806 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 209610 201454
rect 209846 201218 240330 201454
rect 240566 201218 271050 201454
rect 271286 201218 301770 201454
rect 302006 201218 332490 201454
rect 332726 201218 363210 201454
rect 363446 201218 393930 201454
rect 394166 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 209610 201134
rect 209846 200898 240330 201134
rect 240566 200898 271050 201134
rect 271286 200898 301770 201134
rect 302006 200898 332490 201134
rect 332726 200898 363210 201134
rect 363446 200898 393930 201134
rect 394166 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 194250 183454
rect 194486 183218 224970 183454
rect 225206 183218 255690 183454
rect 255926 183218 286410 183454
rect 286646 183218 317130 183454
rect 317366 183218 347850 183454
rect 348086 183218 378570 183454
rect 378806 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 194250 183134
rect 194486 182898 224970 183134
rect 225206 182898 255690 183134
rect 255926 182898 286410 183134
rect 286646 182898 317130 183134
rect 317366 182898 347850 183134
rect 348086 182898 378570 183134
rect 378806 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 209610 165454
rect 209846 165218 240330 165454
rect 240566 165218 271050 165454
rect 271286 165218 301770 165454
rect 302006 165218 332490 165454
rect 332726 165218 363210 165454
rect 363446 165218 393930 165454
rect 394166 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 209610 165134
rect 209846 164898 240330 165134
rect 240566 164898 271050 165134
rect 271286 164898 301770 165134
rect 302006 164898 332490 165134
rect 332726 164898 363210 165134
rect 363446 164898 393930 165134
rect 394166 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 194250 147454
rect 194486 147218 224970 147454
rect 225206 147218 255690 147454
rect 255926 147218 286410 147454
rect 286646 147218 317130 147454
rect 317366 147218 347850 147454
rect 348086 147218 378570 147454
rect 378806 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 194250 147134
rect 194486 146898 224970 147134
rect 225206 146898 255690 147134
rect 255926 146898 286410 147134
rect 286646 146898 317130 147134
rect 317366 146898 347850 147134
rect 348086 146898 378570 147134
rect 378806 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 209610 129454
rect 209846 129218 240330 129454
rect 240566 129218 271050 129454
rect 271286 129218 301770 129454
rect 302006 129218 332490 129454
rect 332726 129218 363210 129454
rect 363446 129218 393930 129454
rect 394166 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 209610 129134
rect 209846 128898 240330 129134
rect 240566 128898 271050 129134
rect 271286 128898 301770 129134
rect 302006 128898 332490 129134
rect 332726 128898 363210 129134
rect 363446 128898 393930 129134
rect 394166 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 34250 111454
rect 34486 111218 64970 111454
rect 65206 111218 95690 111454
rect 95926 111218 126410 111454
rect 126646 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 194250 111454
rect 194486 111218 224970 111454
rect 225206 111218 255690 111454
rect 255926 111218 286410 111454
rect 286646 111218 317130 111454
rect 317366 111218 347850 111454
rect 348086 111218 378570 111454
rect 378806 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 444250 111454
rect 444486 111218 474970 111454
rect 475206 111218 505690 111454
rect 505926 111218 536410 111454
rect 536646 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 34250 111134
rect 34486 110898 64970 111134
rect 65206 110898 95690 111134
rect 95926 110898 126410 111134
rect 126646 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 194250 111134
rect 194486 110898 224970 111134
rect 225206 110898 255690 111134
rect 255926 110898 286410 111134
rect 286646 110898 317130 111134
rect 317366 110898 347850 111134
rect 348086 110898 378570 111134
rect 378806 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 444250 111134
rect 444486 110898 474970 111134
rect 475206 110898 505690 111134
rect 505926 110898 536410 111134
rect 536646 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 49610 93454
rect 49846 93218 80330 93454
rect 80566 93218 111050 93454
rect 111286 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 209610 93454
rect 209846 93218 240330 93454
rect 240566 93218 271050 93454
rect 271286 93218 301770 93454
rect 302006 93218 332490 93454
rect 332726 93218 363210 93454
rect 363446 93218 393930 93454
rect 394166 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 459610 93454
rect 459846 93218 490330 93454
rect 490566 93218 521050 93454
rect 521286 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 49610 93134
rect 49846 92898 80330 93134
rect 80566 92898 111050 93134
rect 111286 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 209610 93134
rect 209846 92898 240330 93134
rect 240566 92898 271050 93134
rect 271286 92898 301770 93134
rect 302006 92898 332490 93134
rect 332726 92898 363210 93134
rect 363446 92898 393930 93134
rect 394166 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 459610 93134
rect 459846 92898 490330 93134
rect 490566 92898 521050 93134
rect 521286 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 34250 75454
rect 34486 75218 64970 75454
rect 65206 75218 95690 75454
rect 95926 75218 126410 75454
rect 126646 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 194250 75454
rect 194486 75218 224970 75454
rect 225206 75218 255690 75454
rect 255926 75218 286410 75454
rect 286646 75218 317130 75454
rect 317366 75218 347850 75454
rect 348086 75218 378570 75454
rect 378806 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 444250 75454
rect 444486 75218 474970 75454
rect 475206 75218 505690 75454
rect 505926 75218 536410 75454
rect 536646 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 34250 75134
rect 34486 74898 64970 75134
rect 65206 74898 95690 75134
rect 95926 74898 126410 75134
rect 126646 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 194250 75134
rect 194486 74898 224970 75134
rect 225206 74898 255690 75134
rect 255926 74898 286410 75134
rect 286646 74898 317130 75134
rect 317366 74898 347850 75134
rect 348086 74898 378570 75134
rect 378806 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 444250 75134
rect 444486 74898 474970 75134
rect 475206 74898 505690 75134
rect 505926 74898 536410 75134
rect 536646 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 49610 57454
rect 49846 57218 80330 57454
rect 80566 57218 111050 57454
rect 111286 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 209610 57454
rect 209846 57218 240330 57454
rect 240566 57218 271050 57454
rect 271286 57218 301770 57454
rect 302006 57218 332490 57454
rect 332726 57218 363210 57454
rect 363446 57218 393930 57454
rect 394166 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 459610 57454
rect 459846 57218 490330 57454
rect 490566 57218 521050 57454
rect 521286 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 49610 57134
rect 49846 56898 80330 57134
rect 80566 56898 111050 57134
rect 111286 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 209610 57134
rect 209846 56898 240330 57134
rect 240566 56898 271050 57134
rect 271286 56898 301770 57134
rect 302006 56898 332490 57134
rect 332726 56898 363210 57134
rect 363446 56898 393930 57134
rect 394166 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 459610 57134
rect 459846 56898 490330 57134
rect 490566 56898 521050 57134
rect 521286 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 34250 39454
rect 34486 39218 64970 39454
rect 65206 39218 95690 39454
rect 95926 39218 126410 39454
rect 126646 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 194250 39454
rect 194486 39218 224970 39454
rect 225206 39218 255690 39454
rect 255926 39218 286410 39454
rect 286646 39218 317130 39454
rect 317366 39218 347850 39454
rect 348086 39218 378570 39454
rect 378806 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 444250 39454
rect 444486 39218 474970 39454
rect 475206 39218 505690 39454
rect 505926 39218 536410 39454
rect 536646 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 34250 39134
rect 34486 38898 64970 39134
rect 65206 38898 95690 39134
rect 95926 38898 126410 39134
rect 126646 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 194250 39134
rect 194486 38898 224970 39134
rect 225206 38898 255690 39134
rect 255926 38898 286410 39134
rect 286646 38898 317130 39134
rect 317366 38898 347850 39134
rect 348086 38898 378570 39134
rect 378806 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 444250 39134
rect 444486 38898 474970 39134
rect 475206 38898 505690 39134
rect 505926 38898 536410 39134
rect 536646 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use Core  core
timestamp 0
transform 1 0 30000 0 1 30000
box 1066 0 100000 100000
use sky130_sram_1kbyte_1rw1r_32x256_8  dmem
timestamp 0
transform 1 0 210000 0 1 300000
box 0 0 95956 79500
use sky130_sram_1kbyte_1rw1r_32x256_8  imem
timestamp 0
transform 1 0 50000 0 1 300000
box 0 0 95956 79500
use Motor_Top  motor
timestamp 0
transform 1 0 440000 0 1 30000
box 0 0 100000 100000
use WB_InterConnect  wb_inter_connect
timestamp 0
transform 1 0 190000 0 1 30000
box 0 0 220000 220000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 132000 74414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 132000 110414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 252000 218414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 252000 254414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 252000 290414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 132000 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 381500 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 381500 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 381500 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 381500 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 381500 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 381500 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 252000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 252000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 252000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 132000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 132000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 132000 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 132000 78134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 132000 114134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 252000 222134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 252000 258134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 252000 294134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 132000 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 381500 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 381500 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 381500 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 381500 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 381500 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 252000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 252000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 252000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 132000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 132000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 132000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 132000 81854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 132000 117854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 252000 225854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 252000 261854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 252000 297854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 132000 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 381500 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 381500 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 252000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 381500 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 381500 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 381500 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 252000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 252000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 252000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 132000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 132000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 132000 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 132000 49574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 132000 85574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 132000 121574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 252000 229574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 252000 265574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 252000 301574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 381500 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 381500 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 381500 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 252000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 381500 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 381500 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 381500 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 252000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 252000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 252000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 132000 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 132000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 132000 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 132000 63854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 132000 99854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 252000 243854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 252000 279854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 381500 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 381500 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 381500 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 252000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 381500 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 381500 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 252000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 252000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 252000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 132000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 132000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 132000 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 132000 67574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 132000 103574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 252000 211574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 252000 247574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 252000 283574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 132000 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 381500 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 381500 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 381500 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 381500 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 381500 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 381500 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 252000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 252000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 252000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 132000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 132000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 132000 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 132000 56414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 132000 92414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 132000 128414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 252000 236414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 252000 272414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 252000 308414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 381500 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 381500 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 381500 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 252000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 381500 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 381500 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 381500 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 252000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 252000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 132000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 132000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 132000 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 132000 60134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 132000 96134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 132000 132134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 252000 240134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 252000 276134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 381500 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 381500 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 381500 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 252000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 381500 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 381500 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 252000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 252000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 252000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 132000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 132000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 132000 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
