magic
tech sky130A
magscale 1 2
timestamp 1647604496
<< obsli1 >>
rect 1104 2159 28888 27761
<< obsm1 >>
rect 1104 2128 28888 27792
<< metal2 >>
rect 18 29200 74 30000
rect 1950 29200 2006 30000
rect 3238 29200 3294 30000
rect 4526 29200 4582 30000
rect 5814 29200 5870 30000
rect 7102 29200 7158 30000
rect 8390 29200 8446 30000
rect 9678 29200 9734 30000
rect 10966 29200 11022 30000
rect 12254 29200 12310 30000
rect 13542 29200 13598 30000
rect 14830 29200 14886 30000
rect 16118 29200 16174 30000
rect 17406 29200 17462 30000
rect 18694 29200 18750 30000
rect 19982 29200 20038 30000
rect 21270 29200 21326 30000
rect 22558 29200 22614 30000
rect 23846 29200 23902 30000
rect 25134 29200 25190 30000
rect 26422 29200 26478 30000
rect 27710 29200 27766 30000
rect 28998 29200 29054 30000
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 10322 0 10378 800
rect 11610 0 11666 800
rect 12898 0 12954 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 19338 0 19394 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 28354 0 28410 800
<< obsm2 >>
rect 1398 29144 1894 29322
rect 2062 29144 3182 29322
rect 3350 29144 4470 29322
rect 4638 29144 5758 29322
rect 5926 29144 7046 29322
rect 7214 29144 8334 29322
rect 8502 29144 9622 29322
rect 9790 29144 10910 29322
rect 11078 29144 12198 29322
rect 12366 29144 13486 29322
rect 13654 29144 14774 29322
rect 14942 29144 16062 29322
rect 16230 29144 17350 29322
rect 17518 29144 18638 29322
rect 18806 29144 19926 29322
rect 20094 29144 21214 29322
rect 21382 29144 22502 29322
rect 22670 29144 23790 29322
rect 23958 29144 25078 29322
rect 25246 29144 26366 29322
rect 26534 29144 27654 29322
rect 27822 29144 28500 29322
rect 1398 856 28500 29144
rect 1418 31 2538 856
rect 2706 31 3826 856
rect 3994 31 5114 856
rect 5282 31 6402 856
rect 6570 31 7690 856
rect 7858 31 8978 856
rect 9146 31 10266 856
rect 10434 31 11554 856
rect 11722 31 12842 856
rect 13010 31 14130 856
rect 14298 31 15418 856
rect 15586 31 16706 856
rect 16874 31 17994 856
rect 18162 31 19282 856
rect 19450 31 20570 856
rect 20738 31 21858 856
rect 22026 31 23146 856
rect 23314 31 24434 856
rect 24602 31 25722 856
rect 25890 31 27010 856
rect 27178 31 28298 856
rect 28466 31 28500 856
<< metal3 >>
rect 0 28568 800 28688
rect 29200 28568 30000 28688
rect 0 27208 800 27328
rect 29200 27208 30000 27328
rect 0 25848 800 25968
rect 29200 25848 30000 25968
rect 0 24488 800 24608
rect 29200 24488 30000 24608
rect 0 23128 800 23248
rect 29200 23128 30000 23248
rect 0 21768 800 21888
rect 29200 21768 30000 21888
rect 0 20408 800 20528
rect 29200 20408 30000 20528
rect 0 19048 800 19168
rect 29200 19048 30000 19168
rect 0 17688 800 17808
rect 29200 17688 30000 17808
rect 0 16328 800 16448
rect 29200 16328 30000 16448
rect 0 14968 800 15088
rect 29200 14968 30000 15088
rect 0 13608 800 13728
rect 29200 13608 30000 13728
rect 0 12248 800 12368
rect 29200 12248 30000 12368
rect 0 10888 800 11008
rect 29200 10888 30000 11008
rect 0 9528 800 9648
rect 29200 9528 30000 9648
rect 0 8168 800 8288
rect 29200 8168 30000 8288
rect 0 6808 800 6928
rect 29200 6808 30000 6928
rect 0 5448 800 5568
rect 29200 5448 30000 5568
rect 0 4088 800 4208
rect 29200 4088 30000 4208
rect 0 2728 800 2848
rect 29200 2728 30000 2848
rect 0 1368 800 1488
rect 29200 1368 30000 1488
rect 29200 8 30000 128
<< obsm3 >>
rect 880 28488 29120 28661
rect 800 27408 29200 28488
rect 880 27128 29120 27408
rect 800 26048 29200 27128
rect 880 25768 29120 26048
rect 800 24688 29200 25768
rect 880 24408 29120 24688
rect 800 23328 29200 24408
rect 880 23048 29120 23328
rect 800 21968 29200 23048
rect 880 21688 29120 21968
rect 800 20608 29200 21688
rect 880 20328 29120 20608
rect 800 19248 29200 20328
rect 880 18968 29120 19248
rect 800 17888 29200 18968
rect 880 17608 29120 17888
rect 800 16528 29200 17608
rect 880 16248 29120 16528
rect 800 15168 29200 16248
rect 880 14888 29120 15168
rect 800 13808 29200 14888
rect 880 13528 29120 13808
rect 800 12448 29200 13528
rect 880 12168 29120 12448
rect 800 11088 29200 12168
rect 880 10808 29120 11088
rect 800 9728 29200 10808
rect 880 9448 29120 9728
rect 800 8368 29200 9448
rect 880 8088 29120 8368
rect 800 7008 29200 8088
rect 880 6728 29120 7008
rect 800 5648 29200 6728
rect 880 5368 29120 5648
rect 800 4288 29200 5368
rect 880 4008 29120 4288
rect 800 2928 29200 4008
rect 880 2648 29120 2928
rect 800 1568 29200 2648
rect 880 1288 29120 1568
rect 800 208 29200 1288
rect 800 35 29120 208
<< metal4 >>
rect 5576 2128 5896 27792
rect 10208 2128 10528 27792
rect 14840 2128 15160 27792
rect 19472 2128 19792 27792
rect 24104 2128 24424 27792
<< obsm4 >>
rect 13491 6835 14760 26349
rect 15240 6835 19392 26349
rect 19872 6835 24024 26349
rect 24504 6835 25701 26349
<< labels >>
rlabel metal3 s 0 14968 800 15088 6 clock
port 1 nsew signal input
rlabel metal3 s 29200 24488 30000 24608 6 io_rxd
port 2 nsew signal input
rlabel metal3 s 29200 5448 30000 5568 6 io_txd
port 3 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 io_uartInt
port 4 nsew signal output
rlabel metal3 s 29200 23128 30000 23248 6 io_uart_select
port 5 nsew signal input
rlabel metal3 s 29200 17688 30000 17808 6 io_wbs_ack_o
port 6 nsew signal output
rlabel metal2 s 13542 29200 13598 30000 6 io_wbs_data_o[0]
port 7 nsew signal output
rlabel metal2 s 12254 29200 12310 30000 6 io_wbs_data_o[10]
port 8 nsew signal output
rlabel metal3 s 29200 10888 30000 11008 6 io_wbs_data_o[11]
port 9 nsew signal output
rlabel metal2 s 1950 29200 2006 30000 6 io_wbs_data_o[12]
port 10 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 io_wbs_data_o[13]
port 11 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 io_wbs_data_o[14]
port 12 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 io_wbs_data_o[15]
port 13 nsew signal output
rlabel metal3 s 29200 21768 30000 21888 6 io_wbs_data_o[16]
port 14 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 io_wbs_data_o[17]
port 15 nsew signal output
rlabel metal3 s 29200 19048 30000 19168 6 io_wbs_data_o[18]
port 16 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 io_wbs_data_o[19]
port 17 nsew signal output
rlabel metal2 s 27710 29200 27766 30000 6 io_wbs_data_o[1]
port 18 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 io_wbs_data_o[20]
port 19 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 io_wbs_data_o[21]
port 20 nsew signal output
rlabel metal2 s 19982 29200 20038 30000 6 io_wbs_data_o[22]
port 21 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 io_wbs_data_o[23]
port 22 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 io_wbs_data_o[24]
port 23 nsew signal output
rlabel metal2 s 18694 29200 18750 30000 6 io_wbs_data_o[25]
port 24 nsew signal output
rlabel metal3 s 29200 20408 30000 20528 6 io_wbs_data_o[26]
port 25 nsew signal output
rlabel metal2 s 5814 29200 5870 30000 6 io_wbs_data_o[27]
port 26 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 io_wbs_data_o[28]
port 27 nsew signal output
rlabel metal3 s 29200 12248 30000 12368 6 io_wbs_data_o[29]
port 28 nsew signal output
rlabel metal2 s 16118 29200 16174 30000 6 io_wbs_data_o[2]
port 29 nsew signal output
rlabel metal3 s 29200 2728 30000 2848 6 io_wbs_data_o[30]
port 30 nsew signal output
rlabel metal2 s 21270 29200 21326 30000 6 io_wbs_data_o[31]
port 31 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 io_wbs_data_o[3]
port 32 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 io_wbs_data_o[4]
port 33 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 io_wbs_data_o[5]
port 34 nsew signal output
rlabel metal2 s 14830 29200 14886 30000 6 io_wbs_data_o[6]
port 35 nsew signal output
rlabel metal3 s 29200 28568 30000 28688 6 io_wbs_data_o[7]
port 36 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 io_wbs_data_o[8]
port 37 nsew signal output
rlabel metal3 s 29200 8 30000 128 6 io_wbs_data_o[9]
port 38 nsew signal output
rlabel metal3 s 29200 9528 30000 9648 6 io_wbs_m2s_addr[0]
port 39 nsew signal input
rlabel metal2 s 18 29200 74 30000 6 io_wbs_m2s_addr[10]
port 40 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 io_wbs_m2s_addr[11]
port 41 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 io_wbs_m2s_addr[12]
port 42 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 io_wbs_m2s_addr[13]
port 43 nsew signal input
rlabel metal3 s 29200 25848 30000 25968 6 io_wbs_m2s_addr[14]
port 44 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 io_wbs_m2s_addr[15]
port 45 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 io_wbs_m2s_addr[1]
port 46 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 io_wbs_m2s_addr[2]
port 47 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 io_wbs_m2s_addr[3]
port 48 nsew signal input
rlabel metal3 s 29200 8168 30000 8288 6 io_wbs_m2s_addr[4]
port 49 nsew signal input
rlabel metal3 s 29200 4088 30000 4208 6 io_wbs_m2s_addr[5]
port 50 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 io_wbs_m2s_addr[6]
port 51 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 io_wbs_m2s_addr[7]
port 52 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 io_wbs_m2s_addr[8]
port 53 nsew signal input
rlabel metal2 s 8390 29200 8446 30000 6 io_wbs_m2s_addr[9]
port 54 nsew signal input
rlabel metal3 s 29200 6808 30000 6928 6 io_wbs_m2s_data[0]
port 55 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 io_wbs_m2s_data[10]
port 56 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 io_wbs_m2s_data[11]
port 57 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 io_wbs_m2s_data[12]
port 58 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 io_wbs_m2s_data[13]
port 59 nsew signal input
rlabel metal2 s 10966 29200 11022 30000 6 io_wbs_m2s_data[14]
port 60 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 io_wbs_m2s_data[15]
port 61 nsew signal input
rlabel metal2 s 18 0 74 800 6 io_wbs_m2s_data[16]
port 62 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 io_wbs_m2s_data[17]
port 63 nsew signal input
rlabel metal2 s 9678 29200 9734 30000 6 io_wbs_m2s_data[18]
port 64 nsew signal input
rlabel metal2 s 17406 29200 17462 30000 6 io_wbs_m2s_data[19]
port 65 nsew signal input
rlabel metal2 s 26422 29200 26478 30000 6 io_wbs_m2s_data[1]
port 66 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 io_wbs_m2s_data[20]
port 67 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 io_wbs_m2s_data[21]
port 68 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 io_wbs_m2s_data[22]
port 69 nsew signal input
rlabel metal2 s 28998 29200 29054 30000 6 io_wbs_m2s_data[23]
port 70 nsew signal input
rlabel metal2 s 22558 29200 22614 30000 6 io_wbs_m2s_data[24]
port 71 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 io_wbs_m2s_data[25]
port 72 nsew signal input
rlabel metal3 s 29200 27208 30000 27328 6 io_wbs_m2s_data[26]
port 73 nsew signal input
rlabel metal3 s 29200 1368 30000 1488 6 io_wbs_m2s_data[27]
port 74 nsew signal input
rlabel metal2 s 4526 29200 4582 30000 6 io_wbs_m2s_data[28]
port 75 nsew signal input
rlabel metal3 s 29200 14968 30000 15088 6 io_wbs_m2s_data[29]
port 76 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 io_wbs_m2s_data[2]
port 77 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 io_wbs_m2s_data[30]
port 78 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 io_wbs_m2s_data[31]
port 79 nsew signal input
rlabel metal3 s 29200 16328 30000 16448 6 io_wbs_m2s_data[3]
port 80 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 io_wbs_m2s_data[4]
port 81 nsew signal input
rlabel metal2 s 25134 29200 25190 30000 6 io_wbs_m2s_data[5]
port 82 nsew signal input
rlabel metal2 s 23846 29200 23902 30000 6 io_wbs_m2s_data[6]
port 83 nsew signal input
rlabel metal2 s 3238 29200 3294 30000 6 io_wbs_m2s_data[7]
port 84 nsew signal input
rlabel metal2 s 7102 29200 7158 30000 6 io_wbs_m2s_data[8]
port 85 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 io_wbs_m2s_data[9]
port 86 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 io_wbs_m2s_stb
port 87 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 io_wbs_m2s_we
port 88 nsew signal input
rlabel metal3 s 29200 13608 30000 13728 6 reset
port 89 nsew signal input
rlabel metal4 s 5576 2128 5896 27792 6 vccd1
port 90 nsew power input
rlabel metal4 s 14840 2128 15160 27792 6 vccd1
port 90 nsew power input
rlabel metal4 s 24104 2128 24424 27792 6 vccd1
port 90 nsew power input
rlabel metal4 s 10208 2128 10528 27792 6 vssd1
port 91 nsew ground input
rlabel metal4 s 19472 2128 19792 27792 6 vssd1
port 91 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2228938
string GDS_FILE /home/em/mpw/UETRV-ECORE/openlane/UART/runs/UART/results/finishing/UART.magic.gds
string GDS_START 423212
<< end >>

